/*
 * World's Smallest Boykisser
 * Author: torbers
 *
 * VGA Example Code
 * Copyright (c) 2024 Tiny Tapeout LTD
 * SPDX-License-Identifier: Apache-2.0
 * Author: Uri Shaked
 */

`default_nettype none

parameter LOGO_SIZE = 128;  // Size of the logo in pixels
parameter DISPLAY_WIDTH = 640;  // VGA display width
parameter DISPLAY_HEIGHT = 480;  // VGA display height

`define COLOR_WHITE 3'd7

module tt_um_torbers_boykisser (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;

  // Configuration
  wire cfg_tile = ui_in[0];

  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  reg [9:0] prev_y;

  hvsync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );

  reg [9:0] logo_left;
  reg [9:0] logo_top;
  reg dir_x;
  reg dir_y;

  wire [2:0] pixel_value;
  reg [2:0] color_index;
  wire [5:0] color;

  wire [9:0] x = pix_x - logo_left;
  wire [9:0] y = pix_y - logo_top;
  wire logo_pixels = cfg_tile || (x[9:7] == 0 && y[9:7] == 0);

  bitmap_rom rom1 (
      .x(x[6:0]),
      .y(y[6:0]),
      .pixel(pixel_value[2:0])
  );

  palette palette_inst (
      .color_index(color_index),
      .rrggbb(color)
  );

  // RGB output logic
  always @(posedge clk) begin
    color_index <= pixel_value;
    if (~rst_n) begin
      R <= 0;
      G <= 0;
      B <= 0;
    end else begin
      R <= 0;
      G <= 0;
      B <= 0;
      if (video_active && logo_pixels) begin
        R <= color[5:4];
        G <= color[3:2];
        B <= color[1:0];
      end
    end
  end

  // Bouncing logic

  always @(posedge clk) begin
    if (~rst_n) begin
      logo_left <= 200;
      logo_top <= 200;
      dir_y <= 0;
      dir_x <= 1;
      color_index <= 0;
    end else begin
      prev_y <= pix_y;
      if (pix_y == 0 && prev_y != pix_y) begin
        logo_left <= logo_left + (dir_x ? 1 : -1);
        logo_top  <= logo_top + (dir_y ? 1 : -1);
        if (logo_left - 1 == 0 && !dir_x) begin
          dir_x <= 1;
          color_index <= color_index + 1;
        end
        if (logo_left + 1 == DISPLAY_WIDTH - LOGO_SIZE && dir_x) begin
          dir_x <= 0;
          color_index <= color_index + 1;
        end
        if (logo_top - 1 == 0 && !dir_y) begin
          dir_y <= 1;
          color_index <= color_index + 1;
        end
        if (logo_top + 1 == DISPLAY_HEIGHT - LOGO_SIZE && dir_y) begin
          dir_y <= 0;
          color_index <= color_index + 1;
        end
      end
    end
  end


endmodule

`default_nettype none

/*
Video sync generator, used to drive a VGA monitor.
Timing from: https://en.wikipedia.org/wiki/Video_Graphics_Array
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
*/

module vga_sync_generator (
    clk,
    reset,
    hsync,
    vsync,
    display_on,
    hpos,
    vpos
);

  input clk;
  input reset;
  output reg hsync, vsync;
  output display_on;
  output reg [9:0] hpos;
  output reg [9:0] vpos;

  // declarations for TV-simulator sync parameters
  // horizontal constants
  parameter H_DISPLAY = 640;  // horizontal display width
  parameter H_BACK = 48;  // horizontal left border (back porch)
  parameter H_FRONT = 16;  // horizontal right border (front porch)
  parameter H_SYNC = 96;  // horizontal sync width
  // vertical constants
  parameter V_DISPLAY = 480;  // vertical display height
  parameter V_TOP = 33;  // vertical top border
  parameter V_BOTTOM = 10;  // vertical bottom border
  parameter V_SYNC = 2;  // vertical sync # lines
  // derived constants
  parameter H_SYNC_START = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START = V_DISPLAY + V_BOTTOM;
  parameter V_SYNC_END = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
  parameter V_MAX = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

  wire hmaxxed = (hpos == H_MAX) || reset;  // set when hpos is maximum
  wire vmaxxed = (vpos == V_MAX) || reset;  // set when vpos is maximum

  // horizontal position counter
  always @(posedge clk) begin
    hsync <= (hpos >= H_SYNC_START && hpos <= H_SYNC_END);
    if (hmaxxed) hpos <= 0;
    else hpos <= hpos + 1;
  end

  // vertical position counter
  always @(posedge clk) begin
    vsync <= (vpos >= V_SYNC_START && vpos <= V_SYNC_END);
    if (hmaxxed)
      if (vmaxxed) vpos <= 0;
      else vpos <= vpos + 1;
  end

  // display_on is set when beam is in "safe" visible frame
  assign display_on = (hpos < H_DISPLAY) && (vpos < V_DISPLAY);

endmodule

// --------------------------------------------------------

module palette (
    input  wire [2:0] color_index,
    output wire [5:0] rrggbb
);

  reg [5:0] palette[7:0];

  initial begin
    palette[0] = 6'b111111;  // blacck
    palette[1] = 6'b110110;  // pink
    palette[2] = 6'b000000;  // green
    palette[3] = 6'b111000;  // orange
    palette[4] = 6'b110011;  // purple
    palette[5] = 6'b011111;  // yellow 
    palette[6] = 6'b110001;  // red
    palette[7] = 6'b111111;  // white
  end

  assign rrggbb = palette[color_index];

endmodule

// --------------------------------------------------------

module bitmap_rom (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire [2:0] pixel
);

// memutommemticmemlly genermemted pixel memory

// Automatically generated pixel memory

reg [7:0] mem_a [0:2047];
initial begin
    mem_a[0] = 8'b00000000;
    mem_a[1] = 8'b00000000;
    mem_a[2] = 8'b00000000;
    mem_a[3] = 8'b00000000;
    mem_a[4] = 8'b00000000;
    mem_a[5] = 8'b00000000;
    mem_a[6] = 8'b00000000;
    mem_a[7] = 8'b00000000;
    mem_a[8] = 8'b00000000;
    mem_a[9] = 8'b00000000;
    mem_a[10] = 8'b00000000;
    mem_a[11] = 8'b00000000;
    mem_a[12] = 8'b00000000;
    mem_a[13] = 8'b00000000;
    mem_a[14] = 8'b00000000;
    mem_a[15] = 8'b00000000;
    mem_a[16] = 8'b00000000;
    mem_a[17] = 8'b00000000;
    mem_a[18] = 8'b00000000;
    mem_a[19] = 8'b00000000;
    mem_a[20] = 8'b00000000;
    mem_a[21] = 8'b00000000;
    mem_a[22] = 8'b00000000;
    mem_a[23] = 8'b00000000;
    mem_a[24] = 8'b00000000;
    mem_a[25] = 8'b00000000;
    mem_a[26] = 8'b00000000;
    mem_a[27] = 8'b00000000;
    mem_a[28] = 8'b00000000;
    mem_a[29] = 8'b00000000;
    mem_a[30] = 8'b00000000;
    mem_a[31] = 8'b00000000;
    mem_a[32] = 8'b00000000;
    mem_a[33] = 8'b00000000;
    mem_a[34] = 8'b00000000;
    mem_a[35] = 8'b00000000;
    mem_a[36] = 8'b00000000;
    mem_a[37] = 8'b00000000;
    mem_a[38] = 8'b00000000;
    mem_a[39] = 8'b00000000;
    mem_a[40] = 8'b00000000;
    mem_a[41] = 8'b00000000;
    mem_a[42] = 8'b00000000;
    mem_a[43] = 8'b00000000;
    mem_a[44] = 8'b00000000;
    mem_a[45] = 8'b00000000;
    mem_a[46] = 8'b00000000;
    mem_a[47] = 8'b00000000;
    mem_a[48] = 8'b00000000;
    mem_a[49] = 8'b00000000;
    mem_a[50] = 8'b00000000;
    mem_a[51] = 8'b00000000;
    mem_a[52] = 8'b00000000;
    mem_a[53] = 8'b00000000;
    mem_a[54] = 8'b00000000;
    mem_a[55] = 8'b00000000;
    mem_a[56] = 8'b00000000;
    mem_a[57] = 8'b00000000;
    mem_a[58] = 8'b00000000;
    mem_a[59] = 8'b00000000;
    mem_a[60] = 8'b00000000;
    mem_a[61] = 8'b00000000;
    mem_a[62] = 8'b00000000;
    mem_a[63] = 8'b00000000;
    mem_a[64] = 8'b00000000;
    mem_a[65] = 8'b00000000;
    mem_a[66] = 8'b00000000;
    mem_a[67] = 8'b00000000;
    mem_a[68] = 8'b00000000;
    mem_a[69] = 8'b00000000;
    mem_a[70] = 8'b00000000;
    mem_a[71] = 8'b00000000;
    mem_a[72] = 8'b00000000;
    mem_a[73] = 8'b00000000;
    mem_a[74] = 8'b00000000;
    mem_a[75] = 8'b00000000;
    mem_a[76] = 8'b00000000;
    mem_a[77] = 8'b00000000;
    mem_a[78] = 8'b00000000;
    mem_a[79] = 8'b00000000;
    mem_a[80] = 8'b00000000;
    mem_a[81] = 8'b00000000;
    mem_a[82] = 8'b00000000;
    mem_a[83] = 8'b00000000;
    mem_a[84] = 8'b00000000;
    mem_a[85] = 8'b00000000;
    mem_a[86] = 8'b00000000;
    mem_a[87] = 8'b00000000;
    mem_a[88] = 8'b00000000;
    mem_a[89] = 8'b00000000;
    mem_a[90] = 8'b00000000;
    mem_a[91] = 8'b00000000;
    mem_a[92] = 8'b00000000;
    mem_a[93] = 8'b00111000;
    mem_a[94] = 8'b00000000;
    mem_a[95] = 8'b00000000;
    mem_a[96] = 8'b00000000;
    mem_a[97] = 8'b00000000;
    mem_a[98] = 8'b00111100;
    mem_a[99] = 8'b00000000;
    mem_a[100] = 8'b00000000;
    mem_a[101] = 8'b00000000;
    mem_a[102] = 8'b00000000;
    mem_a[103] = 8'b00000000;
    mem_a[104] = 8'b00000000;
    mem_a[105] = 8'b00000000;
    mem_a[106] = 8'b00000000;
    mem_a[107] = 8'b00000000;
    mem_a[108] = 8'b00000000;
    mem_a[109] = 8'b00111111;
    mem_a[110] = 8'b00000000;
    mem_a[111] = 8'b00000000;
    mem_a[112] = 8'b00000000;
    mem_a[113] = 8'b00000000;
    mem_a[114] = 8'b11111100;
    mem_a[115] = 8'b00000000;
    mem_a[116] = 8'b00000000;
    mem_a[117] = 8'b00000000;
    mem_a[118] = 8'b00000000;
    mem_a[119] = 8'b00000000;
    mem_a[120] = 8'b00000000;
    mem_a[121] = 8'b00000000;
    mem_a[122] = 8'b00000000;
    mem_a[123] = 8'b00000000;
    mem_a[124] = 8'b11000000;
    mem_a[125] = 8'b00111111;
    mem_a[126] = 8'b00000000;
    mem_a[127] = 8'b00000000;
    mem_a[128] = 8'b00000000;
    mem_a[129] = 8'b00000000;
    mem_a[130] = 8'b11111100;
    mem_a[131] = 8'b00000011;
    mem_a[132] = 8'b00000000;
    mem_a[133] = 8'b00000000;
    mem_a[134] = 8'b00000000;
    mem_a[135] = 8'b00000000;
    mem_a[136] = 8'b00000000;
    mem_a[137] = 8'b00000000;
    mem_a[138] = 8'b00000000;
    mem_a[139] = 8'b00000000;
    mem_a[140] = 8'b11110000;
    mem_a[141] = 8'b01111111;
    mem_a[142] = 8'b00000000;
    mem_a[143] = 8'b00000000;
    mem_a[144] = 8'b00000000;
    mem_a[145] = 8'b00000000;
    mem_a[146] = 8'b11111110;
    mem_a[147] = 8'b00000111;
    mem_a[148] = 8'b00000000;
    mem_a[149] = 8'b00000000;
    mem_a[150] = 8'b00000000;
    mem_a[151] = 8'b00000000;
    mem_a[152] = 8'b00000000;
    mem_a[153] = 8'b00000000;
    mem_a[154] = 8'b00000000;
    mem_a[155] = 8'b00000000;
    mem_a[156] = 8'b11111100;
    mem_a[157] = 8'b01111111;
    mem_a[158] = 8'b00000000;
    mem_a[159] = 8'b00000000;
    mem_a[160] = 8'b00000000;
    mem_a[161] = 8'b00000000;
    mem_a[162] = 8'b11111110;
    mem_a[163] = 8'b00001111;
    mem_a[164] = 8'b00000000;
    mem_a[165] = 8'b00000000;
    mem_a[166] = 8'b00000000;
    mem_a[167] = 8'b00000000;
    mem_a[168] = 8'b00000000;
    mem_a[169] = 8'b00000000;
    mem_a[170] = 8'b00000000;
    mem_a[171] = 8'b00000000;
    mem_a[172] = 8'b11111111;
    mem_a[173] = 8'b01111111;
    mem_a[174] = 8'b00000000;
    mem_a[175] = 8'b00000000;
    mem_a[176] = 8'b00000000;
    mem_a[177] = 8'b00000000;
    mem_a[178] = 8'b11111110;
    mem_a[179] = 8'b00111111;
    mem_a[180] = 8'b00000000;
    mem_a[181] = 8'b00000000;
    mem_a[182] = 8'b00000000;
    mem_a[183] = 8'b00000000;
    mem_a[184] = 8'b00000000;
    mem_a[185] = 8'b00000000;
    mem_a[186] = 8'b00000000;
    mem_a[187] = 8'b11000000;
    mem_a[188] = 8'b11111111;
    mem_a[189] = 8'b11111111;
    mem_a[190] = 8'b00000000;
    mem_a[191] = 8'b00000000;
    mem_a[192] = 8'b00000000;
    mem_a[193] = 8'b00000000;
    mem_a[194] = 8'b11111111;
    mem_a[195] = 8'b01111111;
    mem_a[196] = 8'b00000000;
    mem_a[197] = 8'b00000000;
    mem_a[198] = 8'b00000000;
    mem_a[199] = 8'b00000000;
    mem_a[200] = 8'b00000000;
    mem_a[201] = 8'b00000000;
    mem_a[202] = 8'b00000000;
    mem_a[203] = 8'b11100000;
    mem_a[204] = 8'b11111111;
    mem_a[205] = 8'b11111111;
    mem_a[206] = 8'b00000000;
    mem_a[207] = 8'b00000000;
    mem_a[208] = 8'b00000000;
    mem_a[209] = 8'b00000000;
    mem_a[210] = 8'b11111111;
    mem_a[211] = 8'b11111111;
    mem_a[212] = 8'b00000000;
    mem_a[213] = 8'b00000000;
    mem_a[214] = 8'b11100000;
    mem_a[215] = 8'b00000001;
    mem_a[216] = 8'b00000000;
    mem_a[217] = 8'b00000000;
    mem_a[218] = 8'b00000000;
    mem_a[219] = 8'b11110000;
    mem_a[220] = 8'b11111111;
    mem_a[221] = 8'b11111111;
    mem_a[222] = 8'b00000000;
    mem_a[223] = 8'b00000000;
    mem_a[224] = 8'b00000000;
    mem_a[225] = 8'b00000000;
    mem_a[226] = 8'b11111111;
    mem_a[227] = 8'b11111111;
    mem_a[228] = 8'b00000011;
    mem_a[229] = 8'b00000000;
    mem_a[230] = 8'b11100000;
    mem_a[231] = 8'b00011111;
    mem_a[232] = 8'b00000000;
    mem_a[233] = 8'b00000000;
    mem_a[234] = 8'b00000000;
    mem_a[235] = 8'b11111000;
    mem_a[236] = 8'b11111111;
    mem_a[237] = 8'b11111111;
    mem_a[238] = 8'b00000000;
    mem_a[239] = 8'b00000000;
    mem_a[240] = 8'b00000000;
    mem_a[241] = 8'b00000000;
    mem_a[242] = 8'b11111111;
    mem_a[243] = 8'b11111111;
    mem_a[244] = 8'b00000111;
    mem_a[245] = 8'b00000000;
    mem_a[246] = 8'b11000000;
    mem_a[247] = 8'b11111111;
    mem_a[248] = 8'b00000000;
    mem_a[249] = 8'b00000000;
    mem_a[250] = 8'b00000000;
    mem_a[251] = 8'b11111100;
    mem_a[252] = 8'b11111111;
    mem_a[253] = 8'b11111111;
    mem_a[254] = 8'b00000001;
    mem_a[255] = 8'b00000000;
    mem_a[256] = 8'b00000000;
    mem_a[257] = 8'b00000000;
    mem_a[258] = 8'b11111111;
    mem_a[259] = 8'b11111111;
    mem_a[260] = 8'b00001111;
    mem_a[261] = 8'b00000000;
    mem_a[262] = 8'b11000000;
    mem_a[263] = 8'b11111111;
    mem_a[264] = 8'b00000011;
    mem_a[265] = 8'b00000000;
    mem_a[266] = 8'b00000000;
    mem_a[267] = 8'b11111110;
    mem_a[268] = 8'b11111111;
    mem_a[269] = 8'b11111111;
    mem_a[270] = 8'b00000001;
    mem_a[271] = 8'b00000000;
    mem_a[272] = 8'b00000000;
    mem_a[273] = 8'b10000000;
    mem_a[274] = 8'b11111111;
    mem_a[275] = 8'b11111111;
    mem_a[276] = 8'b00011111;
    mem_a[277] = 8'b00000000;
    mem_a[278] = 8'b10000000;
    mem_a[279] = 8'b11111111;
    mem_a[280] = 8'b00001111;
    mem_a[281] = 8'b00000000;
    mem_a[282] = 8'b10000000;
    mem_a[283] = 8'b11111111;
    mem_a[284] = 8'b11111111;
    mem_a[285] = 8'b11111111;
    mem_a[286] = 8'b00000001;
    mem_a[287] = 8'b00000000;
    mem_a[288] = 8'b00000000;
    mem_a[289] = 8'b10000000;
    mem_a[290] = 8'b11111111;
    mem_a[291] = 8'b11111111;
    mem_a[292] = 8'b00111111;
    mem_a[293] = 8'b00000000;
    mem_a[294] = 8'b10000000;
    mem_a[295] = 8'b11111111;
    mem_a[296] = 8'b00111111;
    mem_a[297] = 8'b00000000;
    mem_a[298] = 8'b10000000;
    mem_a[299] = 8'b11111111;
    mem_a[300] = 8'b11111111;
    mem_a[301] = 8'b11111111;
    mem_a[302] = 8'b00000001;
    mem_a[303] = 8'b00000000;
    mem_a[304] = 8'b00000000;
    mem_a[305] = 8'b10000000;
    mem_a[306] = 8'b11111111;
    mem_a[307] = 8'b11111111;
    mem_a[308] = 8'b01111111;
    mem_a[309] = 8'b00000000;
    mem_a[310] = 8'b00000000;
    mem_a[311] = 8'b11111111;
    mem_a[312] = 8'b11111111;
    mem_a[313] = 8'b00000000;
    mem_a[314] = 8'b11000000;
    mem_a[315] = 8'b11111111;
    mem_a[316] = 8'b11111111;
    mem_a[317] = 8'b11111111;
    mem_a[318] = 8'b00000011;
    mem_a[319] = 8'b00000000;
    mem_a[320] = 8'b00000000;
    mem_a[321] = 8'b10000000;
    mem_a[322] = 8'b11111111;
    mem_a[323] = 8'b11111111;
    mem_a[324] = 8'b11111111;
    mem_a[325] = 8'b00000000;
    mem_a[326] = 8'b00000000;
    mem_a[327] = 8'b11111110;
    mem_a[328] = 8'b11111111;
    mem_a[329] = 8'b00000001;
    mem_a[330] = 8'b11000000;
    mem_a[331] = 8'b11111111;
    mem_a[332] = 8'b11111111;
    mem_a[333] = 8'b11111111;
    mem_a[334] = 8'b00000011;
    mem_a[335] = 8'b00000000;
    mem_a[336] = 8'b00000000;
    mem_a[337] = 8'b10000000;
    mem_a[338] = 8'b11111111;
    mem_a[339] = 8'b11111111;
    mem_a[340] = 8'b11111111;
    mem_a[341] = 8'b00000001;
    mem_a[342] = 8'b00000000;
    mem_a[343] = 8'b11111100;
    mem_a[344] = 8'b11111111;
    mem_a[345] = 8'b00000111;
    mem_a[346] = 8'b11100000;
    mem_a[347] = 8'b11111111;
    mem_a[348] = 8'b11111111;
    mem_a[349] = 8'b11111111;
    mem_a[350] = 8'b00000011;
    mem_a[351] = 8'b00000000;
    mem_a[352] = 8'b00000000;
    mem_a[353] = 8'b11000000;
    mem_a[354] = 8'b11111111;
    mem_a[355] = 8'b11111111;
    mem_a[356] = 8'b11111111;
    mem_a[357] = 8'b00000011;
    mem_a[358] = 8'b00000000;
    mem_a[359] = 8'b11111000;
    mem_a[360] = 8'b11111111;
    mem_a[361] = 8'b00001111;
    mem_a[362] = 8'b11100000;
    mem_a[363] = 8'b11111111;
    mem_a[364] = 8'b11111111;
    mem_a[365] = 8'b11111111;
    mem_a[366] = 8'b00000011;
    mem_a[367] = 8'b00000000;
    mem_a[368] = 8'b00000000;
    mem_a[369] = 8'b11000000;
    mem_a[370] = 8'b11111111;
    mem_a[371] = 8'b11111111;
    mem_a[372] = 8'b11111111;
    mem_a[373] = 8'b00000111;
    mem_a[374] = 8'b00000000;
    mem_a[375] = 8'b11111000;
    mem_a[376] = 8'b11111111;
    mem_a[377] = 8'b00011111;
    mem_a[378] = 8'b11110000;
    mem_a[379] = 8'b11111111;
    mem_a[380] = 8'b11111111;
    mem_a[381] = 8'b11111111;
    mem_a[382] = 8'b00000111;
    mem_a[383] = 8'b00000000;
    mem_a[384] = 8'b00000000;
    mem_a[385] = 8'b11000000;
    mem_a[386] = 8'b11111111;
    mem_a[387] = 8'b11111111;
    mem_a[388] = 8'b11111111;
    mem_a[389] = 8'b00001111;
    mem_a[390] = 8'b00000000;
    mem_a[391] = 8'b11110000;
    mem_a[392] = 8'b11111111;
    mem_a[393] = 8'b00111111;
    mem_a[394] = 8'b11110000;
    mem_a[395] = 8'b11111111;
    mem_a[396] = 8'b11111111;
    mem_a[397] = 8'b11111111;
    mem_a[398] = 8'b00000111;
    mem_a[399] = 8'b00000000;
    mem_a[400] = 8'b00000000;
    mem_a[401] = 8'b11000000;
    mem_a[402] = 8'b11111111;
    mem_a[403] = 8'b11111111;
    mem_a[404] = 8'b11111111;
    mem_a[405] = 8'b00001111;
    mem_a[406] = 8'b00000000;
    mem_a[407] = 8'b11110000;
    mem_a[408] = 8'b11111111;
    mem_a[409] = 8'b01111111;
    mem_a[410] = 8'b11111000;
    mem_a[411] = 8'b11111111;
    mem_a[412] = 8'b11111111;
    mem_a[413] = 8'b11111111;
    mem_a[414] = 8'b00000111;
    mem_a[415] = 8'b00000000;
    mem_a[416] = 8'b00000000;
    mem_a[417] = 8'b11000000;
    mem_a[418] = 8'b11111111;
    mem_a[419] = 8'b11111111;
    mem_a[420] = 8'b11111111;
    mem_a[421] = 8'b00011111;
    mem_a[422] = 8'b00000000;
    mem_a[423] = 8'b11110000;
    mem_a[424] = 8'b11111111;
    mem_a[425] = 8'b11111111;
    mem_a[426] = 8'b11111000;
    mem_a[427] = 8'b11111111;
    mem_a[428] = 8'b11111111;
    mem_a[429] = 8'b11111111;
    mem_a[430] = 8'b00000111;
    mem_a[431] = 8'b00000000;
    mem_a[432] = 8'b00000000;
    mem_a[433] = 8'b11000000;
    mem_a[434] = 8'b11111111;
    mem_a[435] = 8'b11111111;
    mem_a[436] = 8'b11111111;
    mem_a[437] = 8'b00111111;
    mem_a[438] = 8'b00000000;
    mem_a[439] = 8'b11111100;
    mem_a[440] = 8'b11111111;
    mem_a[441] = 8'b11111111;
    mem_a[442] = 8'b11111000;
    mem_a[443] = 8'b11111111;
    mem_a[444] = 8'b11111111;
    mem_a[445] = 8'b11111111;
    mem_a[446] = 8'b00000111;
    mem_a[447] = 8'b00000000;
    mem_a[448] = 8'b00000000;
    mem_a[449] = 8'b11000000;
    mem_a[450] = 8'b11111111;
    mem_a[451] = 8'b11111111;
    mem_a[452] = 8'b11111111;
    mem_a[453] = 8'b11111111;
    mem_a[454] = 8'b11000000;
    mem_a[455] = 8'b11111111;
    mem_a[456] = 8'b11111111;
    mem_a[457] = 8'b11111111;
    mem_a[458] = 8'b11111111;
    mem_a[459] = 8'b11111111;
    mem_a[460] = 8'b11111111;
    mem_a[461] = 8'b11111111;
    mem_a[462] = 8'b00001111;
    mem_a[463] = 8'b00000000;
    mem_a[464] = 8'b00000000;
    mem_a[465] = 8'b11000000;
    mem_a[466] = 8'b11111111;
    mem_a[467] = 8'b11111111;
    mem_a[468] = 8'b11111111;
    mem_a[469] = 8'b01111111;
    mem_a[470] = 8'b11100000;
    mem_a[471] = 8'b11111111;
    mem_a[472] = 8'b11111111;
    mem_a[473] = 8'b11111111;
    mem_a[474] = 8'b11111111;
    mem_a[475] = 8'b11111111;
    mem_a[476] = 8'b11111111;
    mem_a[477] = 8'b11111111;
    mem_a[478] = 8'b00001111;
    mem_a[479] = 8'b00000000;
    mem_a[480] = 8'b00000000;
    mem_a[481] = 8'b11100000;
    mem_a[482] = 8'b11111111;
    mem_a[483] = 8'b11111111;
    mem_a[484] = 8'b11111111;
    mem_a[485] = 8'b00111111;
    mem_a[486] = 8'b11110000;
    mem_a[487] = 8'b11111111;
    mem_a[488] = 8'b11111111;
    mem_a[489] = 8'b11111111;
    mem_a[490] = 8'b11111111;
    mem_a[491] = 8'b11111111;
    mem_a[492] = 8'b11111111;
    mem_a[493] = 8'b11111111;
    mem_a[494] = 8'b00001111;
    mem_a[495] = 8'b00000000;
    mem_a[496] = 8'b00000000;
    mem_a[497] = 8'b11100000;
    mem_a[498] = 8'b11111111;
    mem_a[499] = 8'b11111111;
    mem_a[500] = 8'b11111111;
    mem_a[501] = 8'b00011111;
    mem_a[502] = 8'b11111000;
    mem_a[503] = 8'b11111111;
    mem_a[504] = 8'b11111111;
    mem_a[505] = 8'b11111111;
    mem_a[506] = 8'b11111111;
    mem_a[507] = 8'b11111111;
    mem_a[508] = 8'b11111111;
    mem_a[509] = 8'b11111111;
    mem_a[510] = 8'b00001111;
    mem_a[511] = 8'b00000000;
    mem_a[512] = 8'b00000000;
    mem_a[513] = 8'b11100000;
    mem_a[514] = 8'b11111111;
    mem_a[515] = 8'b11111111;
    mem_a[516] = 8'b11111111;
    mem_a[517] = 8'b00011111;
    mem_a[518] = 8'b00000000;
    mem_a[519] = 8'b11000000;
    mem_a[520] = 8'b11111111;
    mem_a[521] = 8'b11111111;
    mem_a[522] = 8'b11111111;
    mem_a[523] = 8'b11111111;
    mem_a[524] = 8'b11111111;
    mem_a[525] = 8'b11111111;
    mem_a[526] = 8'b00001111;
    mem_a[527] = 8'b00000000;
    mem_a[528] = 8'b00000000;
    mem_a[529] = 8'b11100000;
    mem_a[530] = 8'b11111111;
    mem_a[531] = 8'b11111111;
    mem_a[532] = 8'b11111111;
    mem_a[533] = 8'b00011111;
    mem_a[534] = 8'b00000000;
    mem_a[535] = 8'b00000000;
    mem_a[536] = 8'b11111110;
    mem_a[537] = 8'b11111111;
    mem_a[538] = 8'b11111111;
    mem_a[539] = 8'b11111111;
    mem_a[540] = 8'b11111111;
    mem_a[541] = 8'b11111111;
    mem_a[542] = 8'b00011111;
    mem_a[543] = 8'b00000000;
    mem_a[544] = 8'b00000000;
    mem_a[545] = 8'b11100000;
    mem_a[546] = 8'b11111111;
    mem_a[547] = 8'b11111111;
    mem_a[548] = 8'b11111111;
    mem_a[549] = 8'b00011111;
    mem_a[550] = 8'b00000000;
    mem_a[551] = 8'b00000000;
    mem_a[552] = 8'b11111110;
    mem_a[553] = 8'b11111111;
    mem_a[554] = 8'b11111111;
    mem_a[555] = 8'b11111111;
    mem_a[556] = 8'b11111111;
    mem_a[557] = 8'b11111111;
    mem_a[558] = 8'b00011111;
    mem_a[559] = 8'b00000000;
    mem_a[560] = 8'b00000000;
    mem_a[561] = 8'b11100000;
    mem_a[562] = 8'b11111111;
    mem_a[563] = 8'b11111111;
    mem_a[564] = 8'b11111111;
    mem_a[565] = 8'b11111111;
    mem_a[566] = 8'b11111111;
    mem_a[567] = 8'b00000111;
    mem_a[568] = 8'b11111110;
    mem_a[569] = 8'b11111111;
    mem_a[570] = 8'b11111111;
    mem_a[571] = 8'b11111111;
    mem_a[572] = 8'b11111111;
    mem_a[573] = 8'b11111111;
    mem_a[574] = 8'b00011111;
    mem_a[575] = 8'b00000000;
    mem_a[576] = 8'b00000000;
    mem_a[577] = 8'b11100000;
    mem_a[578] = 8'b11111111;
    mem_a[579] = 8'b11111111;
    mem_a[580] = 8'b11111111;
    mem_a[581] = 8'b11111111;
    mem_a[582] = 8'b11111111;
    mem_a[583] = 8'b11111111;
    mem_a[584] = 8'b11111111;
    mem_a[585] = 8'b11111111;
    mem_a[586] = 8'b11111111;
    mem_a[587] = 8'b11111111;
    mem_a[588] = 8'b11111111;
    mem_a[589] = 8'b11111111;
    mem_a[590] = 8'b00011111;
    mem_a[591] = 8'b00000000;
    mem_a[592] = 8'b00000000;
    mem_a[593] = 8'b11110000;
    mem_a[594] = 8'b11111111;
    mem_a[595] = 8'b11111111;
    mem_a[596] = 8'b11111111;
    mem_a[597] = 8'b11111111;
    mem_a[598] = 8'b11111111;
    mem_a[599] = 8'b11111111;
    mem_a[600] = 8'b11111111;
    mem_a[601] = 8'b11111111;
    mem_a[602] = 8'b11111111;
    mem_a[603] = 8'b11111111;
    mem_a[604] = 8'b11111111;
    mem_a[605] = 8'b11111111;
    mem_a[606] = 8'b00011111;
    mem_a[607] = 8'b00000000;
    mem_a[608] = 8'b00000000;
    mem_a[609] = 8'b11110000;
    mem_a[610] = 8'b11111111;
    mem_a[611] = 8'b11111111;
    mem_a[612] = 8'b11111111;
    mem_a[613] = 8'b11111111;
    mem_a[614] = 8'b11111111;
    mem_a[615] = 8'b11111111;
    mem_a[616] = 8'b11111111;
    mem_a[617] = 8'b11111111;
    mem_a[618] = 8'b11111111;
    mem_a[619] = 8'b11111111;
    mem_a[620] = 8'b11111111;
    mem_a[621] = 8'b11111111;
    mem_a[622] = 8'b00011111;
    mem_a[623] = 8'b00000000;
    mem_a[624] = 8'b00000000;
    mem_a[625] = 8'b11110000;
    mem_a[626] = 8'b11111111;
    mem_a[627] = 8'b11111111;
    mem_a[628] = 8'b11111111;
    mem_a[629] = 8'b11111111;
    mem_a[630] = 8'b11111111;
    mem_a[631] = 8'b11111111;
    mem_a[632] = 8'b11111111;
    mem_a[633] = 8'b11111111;
    mem_a[634] = 8'b11111111;
    mem_a[635] = 8'b11111111;
    mem_a[636] = 8'b11111111;
    mem_a[637] = 8'b11111111;
    mem_a[638] = 8'b00011111;
    mem_a[639] = 8'b00000000;
    mem_a[640] = 8'b00000000;
    mem_a[641] = 8'b11100000;
    mem_a[642] = 8'b11111111;
    mem_a[643] = 8'b11111111;
    mem_a[644] = 8'b11111111;
    mem_a[645] = 8'b11111111;
    mem_a[646] = 8'b11111111;
    mem_a[647] = 8'b11111111;
    mem_a[648] = 8'b11111111;
    mem_a[649] = 8'b11111111;
    mem_a[650] = 8'b11111111;
    mem_a[651] = 8'b11111111;
    mem_a[652] = 8'b11111111;
    mem_a[653] = 8'b11111111;
    mem_a[654] = 8'b00011111;
    mem_a[655] = 8'b00000000;
    mem_a[656] = 8'b00000000;
    mem_a[657] = 8'b11100000;
    mem_a[658] = 8'b11111111;
    mem_a[659] = 8'b11111111;
    mem_a[660] = 8'b11111111;
    mem_a[661] = 8'b11111111;
    mem_a[662] = 8'b11111111;
    mem_a[663] = 8'b11111111;
    mem_a[664] = 8'b11111111;
    mem_a[665] = 8'b11111111;
    mem_a[666] = 8'b11111111;
    mem_a[667] = 8'b11111111;
    mem_a[668] = 8'b11111111;
    mem_a[669] = 8'b11111111;
    mem_a[670] = 8'b00001111;
    mem_a[671] = 8'b00000000;
    mem_a[672] = 8'b00000000;
    mem_a[673] = 8'b11100000;
    mem_a[674] = 8'b11111111;
    mem_a[675] = 8'b11111111;
    mem_a[676] = 8'b11111111;
    mem_a[677] = 8'b11111111;
    mem_a[678] = 8'b11111111;
    mem_a[679] = 8'b11111111;
    mem_a[680] = 8'b11111111;
    mem_a[681] = 8'b11111111;
    mem_a[682] = 8'b11111111;
    mem_a[683] = 8'b11111111;
    mem_a[684] = 8'b11111111;
    mem_a[685] = 8'b11111111;
    mem_a[686] = 8'b00001111;
    mem_a[687] = 8'b00000000;
    mem_a[688] = 8'b00000000;
    mem_a[689] = 8'b11100000;
    mem_a[690] = 8'b11111111;
    mem_a[691] = 8'b11111111;
    mem_a[692] = 8'b11111111;
    mem_a[693] = 8'b11111111;
    mem_a[694] = 8'b11111111;
    mem_a[695] = 8'b11111111;
    mem_a[696] = 8'b11111111;
    mem_a[697] = 8'b11111111;
    mem_a[698] = 8'b11111111;
    mem_a[699] = 8'b11111111;
    mem_a[700] = 8'b11111111;
    mem_a[701] = 8'b11111111;
    mem_a[702] = 8'b00001111;
    mem_a[703] = 8'b00000000;
    mem_a[704] = 8'b00000000;
    mem_a[705] = 8'b11000000;
    mem_a[706] = 8'b11111111;
    mem_a[707] = 8'b11111111;
    mem_a[708] = 8'b11111111;
    mem_a[709] = 8'b11111111;
    mem_a[710] = 8'b11111111;
    mem_a[711] = 8'b11111111;
    mem_a[712] = 8'b11111111;
    mem_a[713] = 8'b11111111;
    mem_a[714] = 8'b11111111;
    mem_a[715] = 8'b11111111;
    mem_a[716] = 8'b11111111;
    mem_a[717] = 8'b11111111;
    mem_a[718] = 8'b00001111;
    mem_a[719] = 8'b00000000;
    mem_a[720] = 8'b00000000;
    mem_a[721] = 8'b11000000;
    mem_a[722] = 8'b11111111;
    mem_a[723] = 8'b11111111;
    mem_a[724] = 8'b11111111;
    mem_a[725] = 8'b11111111;
    mem_a[726] = 8'b11111111;
    mem_a[727] = 8'b11111111;
    mem_a[728] = 8'b11111111;
    mem_a[729] = 8'b11111111;
    mem_a[730] = 8'b11111111;
    mem_a[731] = 8'b11111111;
    mem_a[732] = 8'b11111111;
    mem_a[733] = 8'b11111111;
    mem_a[734] = 8'b00001111;
    mem_a[735] = 8'b00000000;
    mem_a[736] = 8'b00000000;
    mem_a[737] = 8'b11000000;
    mem_a[738] = 8'b11111111;
    mem_a[739] = 8'b11111111;
    mem_a[740] = 8'b11111111;
    mem_a[741] = 8'b11111111;
    mem_a[742] = 8'b11111111;
    mem_a[743] = 8'b11111111;
    mem_a[744] = 8'b11111111;
    mem_a[745] = 8'b11111111;
    mem_a[746] = 8'b11111111;
    mem_a[747] = 8'b11111111;
    mem_a[748] = 8'b11111111;
    mem_a[749] = 8'b11111111;
    mem_a[750] = 8'b00000111;
    mem_a[751] = 8'b00000000;
    mem_a[752] = 8'b00000000;
    mem_a[753] = 8'b10000000;
    mem_a[754] = 8'b11111111;
    mem_a[755] = 8'b11111111;
    mem_a[756] = 8'b11111111;
    mem_a[757] = 8'b11111111;
    mem_a[758] = 8'b11111111;
    mem_a[759] = 8'b11111111;
    mem_a[760] = 8'b11111111;
    mem_a[761] = 8'b11111111;
    mem_a[762] = 8'b11111111;
    mem_a[763] = 8'b11111111;
    mem_a[764] = 8'b11111111;
    mem_a[765] = 8'b11111111;
    mem_a[766] = 8'b00000111;
    mem_a[767] = 8'b00000000;
    mem_a[768] = 8'b00000000;
    mem_a[769] = 8'b10000000;
    mem_a[770] = 8'b11111111;
    mem_a[771] = 8'b11111111;
    mem_a[772] = 8'b11111111;
    mem_a[773] = 8'b11111111;
    mem_a[774] = 8'b11111111;
    mem_a[775] = 8'b11111111;
    mem_a[776] = 8'b11111111;
    mem_a[777] = 8'b11111111;
    mem_a[778] = 8'b11111111;
    mem_a[779] = 8'b11111111;
    mem_a[780] = 8'b11111111;
    mem_a[781] = 8'b11111111;
    mem_a[782] = 8'b00000011;
    mem_a[783] = 8'b00000000;
    mem_a[784] = 8'b00000000;
    mem_a[785] = 8'b00000000;
    mem_a[786] = 8'b11111111;
    mem_a[787] = 8'b11111111;
    mem_a[788] = 8'b11111111;
    mem_a[789] = 8'b11111111;
    mem_a[790] = 8'b11111111;
    mem_a[791] = 8'b11111111;
    mem_a[792] = 8'b11111111;
    mem_a[793] = 8'b11111111;
    mem_a[794] = 8'b11111111;
    mem_a[795] = 8'b11111111;
    mem_a[796] = 8'b11111111;
    mem_a[797] = 8'b11111111;
    mem_a[798] = 8'b00000001;
    mem_a[799] = 8'b00000000;
    mem_a[800] = 8'b00000000;
    mem_a[801] = 8'b00000000;
    mem_a[802] = 8'b11111111;
    mem_a[803] = 8'b11111111;
    mem_a[804] = 8'b11111111;
    mem_a[805] = 8'b11111111;
    mem_a[806] = 8'b11111111;
    mem_a[807] = 8'b11111111;
    mem_a[808] = 8'b11111111;
    mem_a[809] = 8'b01111111;
    mem_a[810] = 8'b00000000;
    mem_a[811] = 8'b00000000;
    mem_a[812] = 8'b11110000;
    mem_a[813] = 8'b11111111;
    mem_a[814] = 8'b00000001;
    mem_a[815] = 8'b00000000;
    mem_a[816] = 8'b00000000;
    mem_a[817] = 8'b00000000;
    mem_a[818] = 8'b11111111;
    mem_a[819] = 8'b11111111;
    mem_a[820] = 8'b11111111;
    mem_a[821] = 8'b11111111;
    mem_a[822] = 8'b11111111;
    mem_a[823] = 8'b11111111;
    mem_a[824] = 8'b11111111;
    mem_a[825] = 8'b00011111;
    mem_a[826] = 8'b00000000;
    mem_a[827] = 8'b00000000;
    mem_a[828] = 8'b11110000;
    mem_a[829] = 8'b11111111;
    mem_a[830] = 8'b00000000;
    mem_a[831] = 8'b00000000;
    mem_a[832] = 8'b00000000;
    mem_a[833] = 8'b00000000;
    mem_a[834] = 8'b11111110;
    mem_a[835] = 8'b00000111;
    mem_a[836] = 8'b00000000;
    mem_a[837] = 8'b00000000;
    mem_a[838] = 8'b11111000;
    mem_a[839] = 8'b11111111;
    mem_a[840] = 8'b11111111;
    mem_a[841] = 8'b00000111;
    mem_a[842] = 8'b00000000;
    mem_a[843] = 8'b00000000;
    mem_a[844] = 8'b11110000;
    mem_a[845] = 8'b01111111;
    mem_a[846] = 8'b00000000;
    mem_a[847] = 8'b00000000;
    mem_a[848] = 8'b00000000;
    mem_a[849] = 8'b00000000;
    mem_a[850] = 8'b11111110;
    mem_a[851] = 8'b00000111;
    mem_a[852] = 8'b00000000;
    mem_a[853] = 8'b00000000;
    mem_a[854] = 8'b11100000;
    mem_a[855] = 8'b11111111;
    mem_a[856] = 8'b11111111;
    mem_a[857] = 8'b00000111;
    mem_a[858] = 8'b10000000;
    mem_a[859] = 8'b00001111;
    mem_a[860] = 8'b11111110;
    mem_a[861] = 8'b00111111;
    mem_a[862] = 8'b00000000;
    mem_a[863] = 8'b00000000;
    mem_a[864] = 8'b00000000;
    mem_a[865] = 8'b00000000;
    mem_a[866] = 8'b11111110;
    mem_a[867] = 8'b00000111;
    mem_a[868] = 8'b00000000;
    mem_a[869] = 8'b00000000;
    mem_a[870] = 8'b11100000;
    mem_a[871] = 8'b11111111;
    mem_a[872] = 8'b11111111;
    mem_a[873] = 8'b00000111;
    mem_a[874] = 8'b10000000;
    mem_a[875] = 8'b00001111;
    mem_a[876] = 8'b11111110;
    mem_a[877] = 8'b00011111;
    mem_a[878] = 8'b00000000;
    mem_a[879] = 8'b00000000;
    mem_a[880] = 8'b00000000;
    mem_a[881] = 8'b00000000;
    mem_a[882] = 8'b11111100;
    mem_a[883] = 8'b00111111;
    mem_a[884] = 8'b11111000;
    mem_a[885] = 8'b00000000;
    mem_a[886] = 8'b11000000;
    mem_a[887] = 8'b11111111;
    mem_a[888] = 8'b11111111;
    mem_a[889] = 8'b00000011;
    mem_a[890] = 8'b10000000;
    mem_a[891] = 8'b00011111;
    mem_a[892] = 8'b11111110;
    mem_a[893] = 8'b00001111;
    mem_a[894] = 8'b00000000;
    mem_a[895] = 8'b00000000;
    mem_a[896] = 8'b00000000;
    mem_a[897] = 8'b00000000;
    mem_a[898] = 8'b11111100;
    mem_a[899] = 8'b00011111;
    mem_a[900] = 8'b11111000;
    mem_a[901] = 8'b00000000;
    mem_a[902] = 8'b11000000;
    mem_a[903] = 8'b11111111;
    mem_a[904] = 8'b11111111;
    mem_a[905] = 8'b00000011;
    mem_a[906] = 8'b10000000;
    mem_a[907] = 8'b00111111;
    mem_a[908] = 8'b11111100;
    mem_a[909] = 8'b00001111;
    mem_a[910] = 8'b00000000;
    mem_a[911] = 8'b00000000;
    mem_a[912] = 8'b00000000;
    mem_a[913] = 8'b00000000;
    mem_a[914] = 8'b11111000;
    mem_a[915] = 8'b00011111;
    mem_a[916] = 8'b11111100;
    mem_a[917] = 8'b00000000;
    mem_a[918] = 8'b11000000;
    mem_a[919] = 8'b11111111;
    mem_a[920] = 8'b11111111;
    mem_a[921] = 8'b00000011;
    mem_a[922] = 8'b10000000;
    mem_a[923] = 8'b00111111;
    mem_a[924] = 8'b11111100;
    mem_a[925] = 8'b00000011;
    mem_a[926] = 8'b00000000;
    mem_a[927] = 8'b00000000;
    mem_a[928] = 8'b00000000;
    mem_a[929] = 8'b00000000;
    mem_a[930] = 8'b11111000;
    mem_a[931] = 8'b00001111;
    mem_a[932] = 8'b11111110;
    mem_a[933] = 8'b00000000;
    mem_a[934] = 8'b11000000;
    mem_a[935] = 8'b11111111;
    mem_a[936] = 8'b11111111;
    mem_a[937] = 8'b00000011;
    mem_a[938] = 8'b10000000;
    mem_a[939] = 8'b01111111;
    mem_a[940] = 8'b11111100;
    mem_a[941] = 8'b00000001;
    mem_a[942] = 8'b00000000;
    mem_a[943] = 8'b00000000;
    mem_a[944] = 8'b00000000;
    mem_a[945] = 8'b00000000;
    mem_a[946] = 8'b11110000;
    mem_a[947] = 8'b00001111;
    mem_a[948] = 8'b11111111;
    mem_a[949] = 8'b00000000;
    mem_a[950] = 8'b11000000;
    mem_a[951] = 8'b11111111;
    mem_a[952] = 8'b11111111;
    mem_a[953] = 8'b00000011;
    mem_a[954] = 8'b10000000;
    mem_a[955] = 8'b01111111;
    mem_a[956] = 8'b11111100;
    mem_a[957] = 8'b00000000;
    mem_a[958] = 8'b00000000;
    mem_a[959] = 8'b00000000;
    mem_a[960] = 8'b00000000;
    mem_a[961] = 8'b00000000;
    mem_a[962] = 8'b11110000;
    mem_a[963] = 8'b00001111;
    mem_a[964] = 8'b11111111;
    mem_a[965] = 8'b00000000;
    mem_a[966] = 8'b11000000;
    mem_a[967] = 8'b11111111;
    mem_a[968] = 8'b11111111;
    mem_a[969] = 8'b00000011;
    mem_a[970] = 8'b10000000;
    mem_a[971] = 8'b01111111;
    mem_a[972] = 8'b11111000;
    mem_a[973] = 8'b00000000;
    mem_a[974] = 8'b00000000;
    mem_a[975] = 8'b00000000;
    mem_a[976] = 8'b00000000;
    mem_a[977] = 8'b00000000;
    mem_a[978] = 8'b11100000;
    mem_a[979] = 8'b10000111;
    mem_a[980] = 8'b11111111;
    mem_a[981] = 8'b00000000;
    mem_a[982] = 8'b11000000;
    mem_a[983] = 8'b11111111;
    mem_a[984] = 8'b11111111;
    mem_a[985] = 8'b00000011;
    mem_a[986] = 8'b10000000;
    mem_a[987] = 8'b01111111;
    mem_a[988] = 8'b11111000;
    mem_a[989] = 8'b00000000;
    mem_a[990] = 8'b00111100;
    mem_a[991] = 8'b00000000;
    mem_a[992] = 8'b00000000;
    mem_a[993] = 8'b00000000;
    mem_a[994] = 8'b11100000;
    mem_a[995] = 8'b10000111;
    mem_a[996] = 8'b11111111;
    mem_a[997] = 8'b00000000;
    mem_a[998] = 8'b11000000;
    mem_a[999] = 8'b11111111;
    mem_a[1000] = 8'b11111111;
    mem_a[1001] = 8'b00000011;
    mem_a[1002] = 8'b10000000;
    mem_a[1003] = 8'b01111111;
    mem_a[1004] = 8'b11111000;
    mem_a[1005] = 8'b11111000;
    mem_a[1006] = 8'b00011111;
    mem_a[1007] = 8'b00000000;
    mem_a[1008] = 8'b00000000;
    mem_a[1009] = 8'b00000000;
    mem_a[1010] = 8'b00000000;
    mem_a[1011] = 8'b10000110;
    mem_a[1012] = 8'b11111111;
    mem_a[1013] = 8'b00000000;
    mem_a[1014] = 8'b11000000;
    mem_a[1015] = 8'b11111111;
    mem_a[1016] = 8'b11111111;
    mem_a[1017] = 8'b00000011;
    mem_a[1018] = 8'b10000000;
    mem_a[1019] = 8'b11111111;
    mem_a[1020] = 8'b11111000;
    mem_a[1021] = 8'b11111111;
    mem_a[1022] = 8'b00011111;
    mem_a[1023] = 8'b00000000;
    mem_a[1024] = 8'b00000000;
    mem_a[1025] = 8'b00000000;
    mem_a[1026] = 8'b00000000;
    mem_a[1027] = 8'b11000110;
    mem_a[1028] = 8'b11111111;
    mem_a[1029] = 8'b00000000;
    mem_a[1030] = 8'b11100000;
    mem_a[1031] = 8'b11111111;
    mem_a[1032] = 8'b11111111;
    mem_a[1033] = 8'b00000011;
    mem_a[1034] = 8'b10000000;
    mem_a[1035] = 8'b11111111;
    mem_a[1036] = 8'b11111000;
    mem_a[1037] = 8'b11111111;
    mem_a[1038] = 8'b00001111;
    mem_a[1039] = 8'b00000000;
    mem_a[1040] = 8'b00000000;
    mem_a[1041] = 8'b00000000;
    mem_a[1042] = 8'b00000000;
    mem_a[1043] = 8'b11000110;
    mem_a[1044] = 8'b11111111;
    mem_a[1045] = 8'b00000000;
    mem_a[1046] = 8'b11100000;
    mem_a[1047] = 8'b11111111;
    mem_a[1048] = 8'b11111111;
    mem_a[1049] = 8'b00000011;
    mem_a[1050] = 8'b10000000;
    mem_a[1051] = 8'b11111111;
    mem_a[1052] = 8'b11111000;
    mem_a[1053] = 8'b11111111;
    mem_a[1054] = 8'b00000111;
    mem_a[1055] = 8'b00000000;
    mem_a[1056] = 8'b00000000;
    mem_a[1057] = 8'b11111000;
    mem_a[1058] = 8'b11111111;
    mem_a[1059] = 8'b11000111;
    mem_a[1060] = 8'b11111111;
    mem_a[1061] = 8'b00000000;
    mem_a[1062] = 8'b11100000;
    mem_a[1063] = 8'b11111111;
    mem_a[1064] = 8'b11111111;
    mem_a[1065] = 8'b00000011;
    mem_a[1066] = 8'b10000000;
    mem_a[1067] = 8'b01111111;
    mem_a[1068] = 8'b11111000;
    mem_a[1069] = 8'b11111111;
    mem_a[1070] = 8'b00000011;
    mem_a[1071] = 8'b00000000;
    mem_a[1072] = 8'b00000000;
    mem_a[1073] = 8'b11110000;
    mem_a[1074] = 8'b11111111;
    mem_a[1075] = 8'b10000111;
    mem_a[1076] = 8'b11111111;
    mem_a[1077] = 8'b00000001;
    mem_a[1078] = 8'b11110000;
    mem_a[1079] = 8'b11111111;
    mem_a[1080] = 8'b11111111;
    mem_a[1081] = 8'b00000111;
    mem_a[1082] = 8'b11000000;
    mem_a[1083] = 8'b01111111;
    mem_a[1084] = 8'b11111000;
    mem_a[1085] = 8'b11111111;
    mem_a[1086] = 8'b00000001;
    mem_a[1087] = 8'b00000000;
    mem_a[1088] = 8'b00000000;
    mem_a[1089] = 8'b11100000;
    mem_a[1090] = 8'b11111111;
    mem_a[1091] = 8'b10000111;
    mem_a[1092] = 8'b11111111;
    mem_a[1093] = 8'b00000001;
    mem_a[1094] = 8'b11110000;
    mem_a[1095] = 8'b11111111;
    mem_a[1096] = 8'b11111111;
    mem_a[1097] = 8'b00000111;
    mem_a[1098] = 8'b11000000;
    mem_a[1099] = 8'b01111111;
    mem_a[1100] = 8'b11111000;
    mem_a[1101] = 8'b01111111;
    mem_a[1102] = 8'b00000000;
    mem_a[1103] = 8'b00000000;
    mem_a[1104] = 8'b00000000;
    mem_a[1105] = 8'b11000000;
    mem_a[1106] = 8'b11111111;
    mem_a[1107] = 8'b10000111;
    mem_a[1108] = 8'b11111111;
    mem_a[1109] = 8'b00000011;
    mem_a[1110] = 8'b11111000;
    mem_a[1111] = 8'b11111111;
    mem_a[1112] = 8'b11111111;
    mem_a[1113] = 8'b00001111;
    mem_a[1114] = 8'b11100000;
    mem_a[1115] = 8'b01111111;
    mem_a[1116] = 8'b11111100;
    mem_a[1117] = 8'b01111111;
    mem_a[1118] = 8'b00000000;
    mem_a[1119] = 8'b00000000;
    mem_a[1120] = 8'b00000000;
    mem_a[1121] = 8'b10000000;
    mem_a[1122] = 8'b11111111;
    mem_a[1123] = 8'b00001111;
    mem_a[1124] = 8'b11111111;
    mem_a[1125] = 8'b00000011;
    mem_a[1126] = 8'b11111100;
    mem_a[1127] = 8'b11111111;
    mem_a[1128] = 8'b11111111;
    mem_a[1129] = 8'b00111111;
    mem_a[1130] = 8'b11111000;
    mem_a[1131] = 8'b01111111;
    mem_a[1132] = 8'b11111100;
    mem_a[1133] = 8'b00111111;
    mem_a[1134] = 8'b00000000;
    mem_a[1135] = 8'b00000000;
    mem_a[1136] = 8'b00000000;
    mem_a[1137] = 8'b00000000;
    mem_a[1138] = 8'b11111111;
    mem_a[1139] = 8'b00001111;
    mem_a[1140] = 8'b11111111;
    mem_a[1141] = 8'b00000111;
    mem_a[1142] = 8'b11111110;
    mem_a[1143] = 8'b11111111;
    mem_a[1144] = 8'b11111111;
    mem_a[1145] = 8'b11111111;
    mem_a[1146] = 8'b11111111;
    mem_a[1147] = 8'b11111111;
    mem_a[1148] = 8'b11111111;
    mem_a[1149] = 8'b00011111;
    mem_a[1150] = 8'b00000000;
    mem_a[1151] = 8'b00000000;
    mem_a[1152] = 8'b00000000;
    mem_a[1153] = 8'b00000000;
    mem_a[1154] = 8'b11111110;
    mem_a[1155] = 8'b00001111;
    mem_a[1156] = 8'b11111111;
    mem_a[1157] = 8'b11111111;
    mem_a[1158] = 8'b11111111;
    mem_a[1159] = 8'b00000000;
    mem_a[1160] = 8'b11111111;
    mem_a[1161] = 8'b11111111;
    mem_a[1162] = 8'b11111111;
    mem_a[1163] = 8'b11111111;
    mem_a[1164] = 8'b11111111;
    mem_a[1165] = 8'b00001111;
    mem_a[1166] = 8'b00000000;
    mem_a[1167] = 8'b00000000;
    mem_a[1168] = 8'b00000000;
    mem_a[1169] = 8'b00000000;
    mem_a[1170] = 8'b11111100;
    mem_a[1171] = 8'b00011111;
    mem_a[1172] = 8'b11111111;
    mem_a[1173] = 8'b11111111;
    mem_a[1174] = 8'b11111111;
    mem_a[1175] = 8'b00000000;
    mem_a[1176] = 8'b11111111;
    mem_a[1177] = 8'b11111111;
    mem_a[1178] = 8'b11111111;
    mem_a[1179] = 8'b11111111;
    mem_a[1180] = 8'b11111111;
    mem_a[1181] = 8'b00001111;
    mem_a[1182] = 8'b00000000;
    mem_a[1183] = 8'b00000000;
    mem_a[1184] = 8'b00000000;
    mem_a[1185] = 8'b00000000;
    mem_a[1186] = 8'b11111000;
    mem_a[1187] = 8'b11111111;
    mem_a[1188] = 8'b11111111;
    mem_a[1189] = 8'b11111111;
    mem_a[1190] = 8'b11111111;
    mem_a[1191] = 8'b00000000;
    mem_a[1192] = 8'b11111111;
    mem_a[1193] = 8'b11111111;
    mem_a[1194] = 8'b11111111;
    mem_a[1195] = 8'b11111111;
    mem_a[1196] = 8'b11111111;
    mem_a[1197] = 8'b00001111;
    mem_a[1198] = 8'b00000000;
    mem_a[1199] = 8'b00000000;
    mem_a[1200] = 8'b00000000;
    mem_a[1201] = 8'b00000000;
    mem_a[1202] = 8'b11111000;
    mem_a[1203] = 8'b11111111;
    mem_a[1204] = 8'b11111111;
    mem_a[1205] = 8'b11111111;
    mem_a[1206] = 8'b11111111;
    mem_a[1207] = 8'b11111111;
    mem_a[1208] = 8'b11111111;
    mem_a[1209] = 8'b11111111;
    mem_a[1210] = 8'b11111111;
    mem_a[1211] = 8'b11111111;
    mem_a[1212] = 8'b11111111;
    mem_a[1213] = 8'b00001111;
    mem_a[1214] = 8'b00000000;
    mem_a[1215] = 8'b00000000;
    mem_a[1216] = 8'b00000000;
    mem_a[1217] = 8'b00000000;
    mem_a[1218] = 8'b11111000;
    mem_a[1219] = 8'b11111111;
    mem_a[1220] = 8'b11111111;
    mem_a[1221] = 8'b11111111;
    mem_a[1222] = 8'b11111111;
    mem_a[1223] = 8'b11111111;
    mem_a[1224] = 8'b11111111;
    mem_a[1225] = 8'b11111111;
    mem_a[1226] = 8'b11111111;
    mem_a[1227] = 8'b11111111;
    mem_a[1228] = 8'b11111111;
    mem_a[1229] = 8'b00011111;
    mem_a[1230] = 8'b00000000;
    mem_a[1231] = 8'b00000000;
    mem_a[1232] = 8'b00000000;
    mem_a[1233] = 8'b00000000;
    mem_a[1234] = 8'b11111000;
    mem_a[1235] = 8'b11111111;
    mem_a[1236] = 8'b11111111;
    mem_a[1237] = 8'b11111111;
    mem_a[1238] = 8'b11111111;
    mem_a[1239] = 8'b11111111;
    mem_a[1240] = 8'b11111111;
    mem_a[1241] = 8'b11111111;
    mem_a[1242] = 8'b11111111;
    mem_a[1243] = 8'b11111111;
    mem_a[1244] = 8'b11111111;
    mem_a[1245] = 8'b00111111;
    mem_a[1246] = 8'b00000000;
    mem_a[1247] = 8'b00000000;
    mem_a[1248] = 8'b00000000;
    mem_a[1249] = 8'b00000000;
    mem_a[1250] = 8'b11111100;
    mem_a[1251] = 8'b11111111;
    mem_a[1252] = 8'b11111111;
    mem_a[1253] = 8'b11111111;
    mem_a[1254] = 8'b11111111;
    mem_a[1255] = 8'b11111111;
    mem_a[1256] = 8'b11111111;
    mem_a[1257] = 8'b11111111;
    mem_a[1258] = 8'b11111111;
    mem_a[1259] = 8'b11111111;
    mem_a[1260] = 8'b11111111;
    mem_a[1261] = 8'b01111111;
    mem_a[1262] = 8'b00000000;
    mem_a[1263] = 8'b00000000;
    mem_a[1264] = 8'b00000000;
    mem_a[1265] = 8'b00000000;
    mem_a[1266] = 8'b11111100;
    mem_a[1267] = 8'b11111111;
    mem_a[1268] = 8'b11111111;
    mem_a[1269] = 8'b11111111;
    mem_a[1270] = 8'b11111111;
    mem_a[1271] = 8'b11111111;
    mem_a[1272] = 8'b11111111;
    mem_a[1273] = 8'b11100011;
    mem_a[1274] = 8'b11111111;
    mem_a[1275] = 8'b11111111;
    mem_a[1276] = 8'b11111111;
    mem_a[1277] = 8'b11111111;
    mem_a[1278] = 8'b00000000;
    mem_a[1279] = 8'b00000000;
    mem_a[1280] = 8'b00000000;
    mem_a[1281] = 8'b00000000;
    mem_a[1282] = 8'b11111110;
    mem_a[1283] = 8'b11111111;
    mem_a[1284] = 8'b11111111;
    mem_a[1285] = 8'b11111111;
    mem_a[1286] = 8'b11111111;
    mem_a[1287] = 8'b00011111;
    mem_a[1288] = 8'b11111111;
    mem_a[1289] = 8'b11100000;
    mem_a[1290] = 8'b11111111;
    mem_a[1291] = 8'b11111111;
    mem_a[1292] = 8'b11111111;
    mem_a[1293] = 8'b11111111;
    mem_a[1294] = 8'b00000001;
    mem_a[1295] = 8'b00000000;
    mem_a[1296] = 8'b00000000;
    mem_a[1297] = 8'b00000000;
    mem_a[1298] = 8'b11111110;
    mem_a[1299] = 8'b11111111;
    mem_a[1300] = 8'b11111111;
    mem_a[1301] = 8'b11111111;
    mem_a[1302] = 8'b11111111;
    mem_a[1303] = 8'b00001111;
    mem_a[1304] = 8'b01111110;
    mem_a[1305] = 8'b11100000;
    mem_a[1306] = 8'b11111111;
    mem_a[1307] = 8'b11111111;
    mem_a[1308] = 8'b11111111;
    mem_a[1309] = 8'b11111111;
    mem_a[1310] = 8'b00000001;
    mem_a[1311] = 8'b00000000;
    mem_a[1312] = 8'b00000000;
    mem_a[1313] = 8'b00000000;
    mem_a[1314] = 8'b11111111;
    mem_a[1315] = 8'b11111111;
    mem_a[1316] = 8'b11111111;
    mem_a[1317] = 8'b11111111;
    mem_a[1318] = 8'b11111111;
    mem_a[1319] = 8'b00000111;
    mem_a[1320] = 8'b00000000;
    mem_a[1321] = 8'b11100000;
    mem_a[1322] = 8'b11111111;
    mem_a[1323] = 8'b11111111;
    mem_a[1324] = 8'b11111111;
    mem_a[1325] = 8'b11111111;
    mem_a[1326] = 8'b00000011;
    mem_a[1327] = 8'b00000000;
    mem_a[1328] = 8'b00000000;
    mem_a[1329] = 8'b00000000;
    mem_a[1330] = 8'b11111111;
    mem_a[1331] = 8'b11111111;
    mem_a[1332] = 8'b11111111;
    mem_a[1333] = 8'b11111111;
    mem_a[1334] = 8'b10000011;
    mem_a[1335] = 8'b00000001;
    mem_a[1336] = 8'b00000000;
    mem_a[1337] = 8'b11111000;
    mem_a[1338] = 8'b11111111;
    mem_a[1339] = 8'b11111111;
    mem_a[1340] = 8'b11111111;
    mem_a[1341] = 8'b11111111;
    mem_a[1342] = 8'b00000011;
    mem_a[1343] = 8'b00000000;
    mem_a[1344] = 8'b00000000;
    mem_a[1345] = 8'b10000000;
    mem_a[1346] = 8'b11111111;
    mem_a[1347] = 8'b11111111;
    mem_a[1348] = 8'b11111111;
    mem_a[1349] = 8'b11111111;
    mem_a[1350] = 8'b00000011;
    mem_a[1351] = 8'b00000000;
    mem_a[1352] = 8'b00000000;
    mem_a[1353] = 8'b11111100;
    mem_a[1354] = 8'b11111111;
    mem_a[1355] = 8'b11111111;
    mem_a[1356] = 8'b11111111;
    mem_a[1357] = 8'b11111111;
    mem_a[1358] = 8'b00000000;
    mem_a[1359] = 8'b00000000;
    mem_a[1360] = 8'b00000000;
    mem_a[1361] = 8'b10000000;
    mem_a[1362] = 8'b11111111;
    mem_a[1363] = 8'b11111111;
    mem_a[1364] = 8'b11111111;
    mem_a[1365] = 8'b11111111;
    mem_a[1366] = 8'b00000011;
    mem_a[1367] = 8'b11000000;
    mem_a[1368] = 8'b10000001;
    mem_a[1369] = 8'b11111111;
    mem_a[1370] = 8'b11111111;
    mem_a[1371] = 8'b11111111;
    mem_a[1372] = 8'b11110000;
    mem_a[1373] = 8'b00111111;
    mem_a[1374] = 8'b00000000;
    mem_a[1375] = 8'b00000000;
    mem_a[1376] = 8'b00000000;
    mem_a[1377] = 8'b10000000;
    mem_a[1378] = 8'b11111111;
    mem_a[1379] = 8'b11111111;
    mem_a[1380] = 8'b11111111;
    mem_a[1381] = 8'b11111111;
    mem_a[1382] = 8'b00001111;
    mem_a[1383] = 8'b11110000;
    mem_a[1384] = 8'b11111111;
    mem_a[1385] = 8'b11111111;
    mem_a[1386] = 8'b11111111;
    mem_a[1387] = 8'b01111111;
    mem_a[1388] = 8'b11110000;
    mem_a[1389] = 8'b00000000;
    mem_a[1390] = 8'b00000000;
    mem_a[1391] = 8'b00000000;
    mem_a[1392] = 8'b00000000;
    mem_a[1393] = 8'b00000000;
    mem_a[1394] = 8'b01111100;
    mem_a[1395] = 8'b10000000;
    mem_a[1396] = 8'b11111111;
    mem_a[1397] = 8'b11111111;
    mem_a[1398] = 8'b11111111;
    mem_a[1399] = 8'b11111111;
    mem_a[1400] = 8'b11111111;
    mem_a[1401] = 8'b11111111;
    mem_a[1402] = 8'b11111111;
    mem_a[1403] = 8'b00111111;
    mem_a[1404] = 8'b00000000;
    mem_a[1405] = 8'b00000000;
    mem_a[1406] = 8'b00000000;
    mem_a[1407] = 8'b00000000;
    mem_a[1408] = 8'b00000000;
    mem_a[1409] = 8'b00000000;
    mem_a[1410] = 8'b00000000;
    mem_a[1411] = 8'b00000000;
    mem_a[1412] = 8'b11111110;
    mem_a[1413] = 8'b11111111;
    mem_a[1414] = 8'b11111111;
    mem_a[1415] = 8'b11111111;
    mem_a[1416] = 8'b11111111;
    mem_a[1417] = 8'b11111111;
    mem_a[1418] = 8'b11111111;
    mem_a[1419] = 8'b00001111;
    mem_a[1420] = 8'b00000000;
    mem_a[1421] = 8'b00000000;
    mem_a[1422] = 8'b00000000;
    mem_a[1423] = 8'b00000000;
    mem_a[1424] = 8'b00000000;
    mem_a[1425] = 8'b00000000;
    mem_a[1426] = 8'b00000000;
    mem_a[1427] = 8'b00000000;
    mem_a[1428] = 8'b11111100;
    mem_a[1429] = 8'b11111111;
    mem_a[1430] = 8'b11111111;
    mem_a[1431] = 8'b11111111;
    mem_a[1432] = 8'b11111111;
    mem_a[1433] = 8'b11111111;
    mem_a[1434] = 8'b11111111;
    mem_a[1435] = 8'b00000011;
    mem_a[1436] = 8'b00000000;
    mem_a[1437] = 8'b00000000;
    mem_a[1438] = 8'b00000000;
    mem_a[1439] = 8'b00000000;
    mem_a[1440] = 8'b00000000;
    mem_a[1441] = 8'b00000000;
    mem_a[1442] = 8'b00000000;
    mem_a[1443] = 8'b00000000;
    mem_a[1444] = 8'b11110000;
    mem_a[1445] = 8'b11111111;
    mem_a[1446] = 8'b11111111;
    mem_a[1447] = 8'b11111111;
    mem_a[1448] = 8'b11111111;
    mem_a[1449] = 8'b11111111;
    mem_a[1450] = 8'b11111111;
    mem_a[1451] = 8'b00000000;
    mem_a[1452] = 8'b00000000;
    mem_a[1453] = 8'b00000000;
    mem_a[1454] = 8'b00000000;
    mem_a[1455] = 8'b00000000;
    mem_a[1456] = 8'b00000000;
    mem_a[1457] = 8'b00000000;
    mem_a[1458] = 8'b00000000;
    mem_a[1459] = 8'b00000000;
    mem_a[1460] = 8'b11000000;
    mem_a[1461] = 8'b11111111;
    mem_a[1462] = 8'b11111111;
    mem_a[1463] = 8'b11111111;
    mem_a[1464] = 8'b11111111;
    mem_a[1465] = 8'b11111111;
    mem_a[1466] = 8'b00011111;
    mem_a[1467] = 8'b00000000;
    mem_a[1468] = 8'b00000000;
    mem_a[1469] = 8'b00000000;
    mem_a[1470] = 8'b00000000;
    mem_a[1471] = 8'b00000000;
    mem_a[1472] = 8'b00000000;
    mem_a[1473] = 8'b00000000;
    mem_a[1474] = 8'b00000000;
    mem_a[1475] = 8'b00000000;
    mem_a[1476] = 8'b00000000;
    mem_a[1477] = 8'b11000000;
    mem_a[1478] = 8'b11111111;
    mem_a[1479] = 8'b11111111;
    mem_a[1480] = 8'b11111111;
    mem_a[1481] = 8'b11111111;
    mem_a[1482] = 8'b00000011;
    mem_a[1483] = 8'b00000000;
    mem_a[1484] = 8'b00000000;
    mem_a[1485] = 8'b00000000;
    mem_a[1486] = 8'b00000000;
    mem_a[1487] = 8'b00000000;
    mem_a[1488] = 8'b00000000;
    mem_a[1489] = 8'b00000000;
    mem_a[1490] = 8'b00000000;
    mem_a[1491] = 8'b00000000;
    mem_a[1492] = 8'b00000000;
    mem_a[1493] = 8'b00000000;
    mem_a[1494] = 8'b11111111;
    mem_a[1495] = 8'b11111111;
    mem_a[1496] = 8'b11111111;
    mem_a[1497] = 8'b11111111;
    mem_a[1498] = 8'b00000011;
    mem_a[1499] = 8'b00000000;
    mem_a[1500] = 8'b00000000;
    mem_a[1501] = 8'b00000000;
    mem_a[1502] = 8'b00000000;
    mem_a[1503] = 8'b00000000;
    mem_a[1504] = 8'b00000000;
    mem_a[1505] = 8'b00000000;
    mem_a[1506] = 8'b00000000;
    mem_a[1507] = 8'b00000000;
    mem_a[1508] = 8'b00000000;
    mem_a[1509] = 8'b00000000;
    mem_a[1510] = 8'b11000000;
    mem_a[1511] = 8'b11111111;
    mem_a[1512] = 8'b11111111;
    mem_a[1513] = 8'b11111111;
    mem_a[1514] = 8'b10000011;
    mem_a[1515] = 8'b00000001;
    mem_a[1516] = 8'b00000000;
    mem_a[1517] = 8'b00000000;
    mem_a[1518] = 8'b00000000;
    mem_a[1519] = 8'b00000000;
    mem_a[1520] = 8'b00000000;
    mem_a[1521] = 8'b00000000;
    mem_a[1522] = 8'b00000000;
    mem_a[1523] = 8'b00000000;
    mem_a[1524] = 8'b00000000;
    mem_a[1525] = 8'b00000110;
    mem_a[1526] = 8'b11000000;
    mem_a[1527] = 8'b11111111;
    mem_a[1528] = 8'b11111111;
    mem_a[1529] = 8'b11111111;
    mem_a[1530] = 8'b11111111;
    mem_a[1531] = 8'b00000001;
    mem_a[1532] = 8'b00000000;
    mem_a[1533] = 8'b00000000;
    mem_a[1534] = 8'b00000000;
    mem_a[1535] = 8'b00000000;
    mem_a[1536] = 8'b00000000;
    mem_a[1537] = 8'b00000000;
    mem_a[1538] = 8'b00000000;
    mem_a[1539] = 8'b00000000;
    mem_a[1540] = 8'b00000000;
    mem_a[1541] = 8'b00111100;
    mem_a[1542] = 8'b11000000;
    mem_a[1543] = 8'b11111111;
    mem_a[1544] = 8'b11111111;
    mem_a[1545] = 8'b11111111;
    mem_a[1546] = 8'b00111111;
    mem_a[1547] = 8'b00000000;
    mem_a[1548] = 8'b00000000;
    mem_a[1549] = 8'b00000000;
    mem_a[1550] = 8'b00000000;
    mem_a[1551] = 8'b00000000;
    mem_a[1552] = 8'b00000000;
    mem_a[1553] = 8'b00000000;
    mem_a[1554] = 8'b00000000;
    mem_a[1555] = 8'b00000000;
    mem_a[1556] = 8'b00000000;
    mem_a[1557] = 8'b11111100;
    mem_a[1558] = 8'b11111111;
    mem_a[1559] = 8'b11111111;
    mem_a[1560] = 8'b11111111;
    mem_a[1561] = 8'b11111111;
    mem_a[1562] = 8'b00111111;
    mem_a[1563] = 8'b00000000;
    mem_a[1564] = 8'b00000000;
    mem_a[1565] = 8'b00000000;
    mem_a[1566] = 8'b00000000;
    mem_a[1567] = 8'b00000000;
    mem_a[1568] = 8'b00000000;
    mem_a[1569] = 8'b00000000;
    mem_a[1570] = 8'b00000000;
    mem_a[1571] = 8'b00000000;
    mem_a[1572] = 8'b00000000;
    mem_a[1573] = 8'b11111000;
    mem_a[1574] = 8'b11111111;
    mem_a[1575] = 8'b11111111;
    mem_a[1576] = 8'b11111111;
    mem_a[1577] = 8'b11111111;
    mem_a[1578] = 8'b00111111;
    mem_a[1579] = 8'b00000000;
    mem_a[1580] = 8'b00000000;
    mem_a[1581] = 8'b00000000;
    mem_a[1582] = 8'b00000000;
    mem_a[1583] = 8'b00000000;
    mem_a[1584] = 8'b00000000;
    mem_a[1585] = 8'b00000000;
    mem_a[1586] = 8'b00000000;
    mem_a[1587] = 8'b00000000;
    mem_a[1588] = 8'b00000000;
    mem_a[1589] = 8'b11110000;
    mem_a[1590] = 8'b11111111;
    mem_a[1591] = 8'b11111111;
    mem_a[1592] = 8'b11111111;
    mem_a[1593] = 8'b11111111;
    mem_a[1594] = 8'b01111111;
    mem_a[1595] = 8'b00000000;
    mem_a[1596] = 8'b00000000;
    mem_a[1597] = 8'b00000000;
    mem_a[1598] = 8'b00000000;
    mem_a[1599] = 8'b00000000;
    mem_a[1600] = 8'b00000000;
    mem_a[1601] = 8'b00000000;
    mem_a[1602] = 8'b00000000;
    mem_a[1603] = 8'b00000000;
    mem_a[1604] = 8'b00000000;
    mem_a[1605] = 8'b11100000;
    mem_a[1606] = 8'b11111111;
    mem_a[1607] = 8'b11111111;
    mem_a[1608] = 8'b11111111;
    mem_a[1609] = 8'b11111111;
    mem_a[1610] = 8'b01111111;
    mem_a[1611] = 8'b00000000;
    mem_a[1612] = 8'b00000000;
    mem_a[1613] = 8'b00000000;
    mem_a[1614] = 8'b00000000;
    mem_a[1615] = 8'b00000000;
    mem_a[1616] = 8'b00000000;
    mem_a[1617] = 8'b00000000;
    mem_a[1618] = 8'b00000000;
    mem_a[1619] = 8'b00000000;
    mem_a[1620] = 8'b00000000;
    mem_a[1621] = 8'b11000000;
    mem_a[1622] = 8'b11111111;
    mem_a[1623] = 8'b11111111;
    mem_a[1624] = 8'b11111111;
    mem_a[1625] = 8'b11111111;
    mem_a[1626] = 8'b11111111;
    mem_a[1627] = 8'b00000000;
    mem_a[1628] = 8'b00000000;
    mem_a[1629] = 8'b00000000;
    mem_a[1630] = 8'b00000000;
    mem_a[1631] = 8'b00000000;
    mem_a[1632] = 8'b00000000;
    mem_a[1633] = 8'b00000000;
    mem_a[1634] = 8'b00000000;
    mem_a[1635] = 8'b00000000;
    mem_a[1636] = 8'b00000000;
    mem_a[1637] = 8'b10000000;
    mem_a[1638] = 8'b11111111;
    mem_a[1639] = 8'b11111111;
    mem_a[1640] = 8'b11111111;
    mem_a[1641] = 8'b11111111;
    mem_a[1642] = 8'b11111111;
    mem_a[1643] = 8'b00000001;
    mem_a[1644] = 8'b00000000;
    mem_a[1645] = 8'b00000000;
    mem_a[1646] = 8'b00000000;
    mem_a[1647] = 8'b00000000;
    mem_a[1648] = 8'b00000000;
    mem_a[1649] = 8'b00000000;
    mem_a[1650] = 8'b00000000;
    mem_a[1651] = 8'b00000000;
    mem_a[1652] = 8'b00000000;
    mem_a[1653] = 8'b10000000;
    mem_a[1654] = 8'b11111111;
    mem_a[1655] = 8'b11111111;
    mem_a[1656] = 8'b11111111;
    mem_a[1657] = 8'b11111111;
    mem_a[1658] = 8'b11111111;
    mem_a[1659] = 8'b00000001;
    mem_a[1660] = 8'b00000000;
    mem_a[1661] = 8'b00000000;
    mem_a[1662] = 8'b00000000;
    mem_a[1663] = 8'b00000000;
    mem_a[1664] = 8'b00000000;
    mem_a[1665] = 8'b00000000;
    mem_a[1666] = 8'b00000000;
    mem_a[1667] = 8'b00000000;
    mem_a[1668] = 8'b00000000;
    mem_a[1669] = 8'b10000000;
    mem_a[1670] = 8'b11111111;
    mem_a[1671] = 8'b11111111;
    mem_a[1672] = 8'b11111111;
    mem_a[1673] = 8'b11111111;
    mem_a[1674] = 8'b11111111;
    mem_a[1675] = 8'b00000011;
    mem_a[1676] = 8'b00000000;
    mem_a[1677] = 8'b00000000;
    mem_a[1678] = 8'b00000000;
    mem_a[1679] = 8'b00000000;
    mem_a[1680] = 8'b00000000;
    mem_a[1681] = 8'b00000000;
    mem_a[1682] = 8'b00000000;
    mem_a[1683] = 8'b00000000;
    mem_a[1684] = 8'b00000000;
    mem_a[1685] = 8'b10000000;
    mem_a[1686] = 8'b11111111;
    mem_a[1687] = 8'b11111111;
    mem_a[1688] = 8'b11111111;
    mem_a[1689] = 8'b11111111;
    mem_a[1690] = 8'b11111111;
    mem_a[1691] = 8'b00000011;
    mem_a[1692] = 8'b00000000;
    mem_a[1693] = 8'b00000000;
    mem_a[1694] = 8'b00000000;
    mem_a[1695] = 8'b00000000;
    mem_a[1696] = 8'b00000000;
    mem_a[1697] = 8'b00000000;
    mem_a[1698] = 8'b00000000;
    mem_a[1699] = 8'b00000000;
    mem_a[1700] = 8'b00000000;
    mem_a[1701] = 8'b10000000;
    mem_a[1702] = 8'b11111111;
    mem_a[1703] = 8'b11111111;
    mem_a[1704] = 8'b11111111;
    mem_a[1705] = 8'b11111111;
    mem_a[1706] = 8'b11111111;
    mem_a[1707] = 8'b00000011;
    mem_a[1708] = 8'b00000000;
    mem_a[1709] = 8'b00000000;
    mem_a[1710] = 8'b00000000;
    mem_a[1711] = 8'b00000000;
    mem_a[1712] = 8'b00000000;
    mem_a[1713] = 8'b00000000;
    mem_a[1714] = 8'b00000000;
    mem_a[1715] = 8'b00000000;
    mem_a[1716] = 8'b00000000;
    mem_a[1717] = 8'b11000000;
    mem_a[1718] = 8'b11111111;
    mem_a[1719] = 8'b11111111;
    mem_a[1720] = 8'b11111111;
    mem_a[1721] = 8'b11111111;
    mem_a[1722] = 8'b11111111;
    mem_a[1723] = 8'b00000111;
    mem_a[1724] = 8'b00000000;
    mem_a[1725] = 8'b00000000;
    mem_a[1726] = 8'b00000000;
    mem_a[1727] = 8'b00000000;
    mem_a[1728] = 8'b00000000;
    mem_a[1729] = 8'b00000000;
    mem_a[1730] = 8'b00000000;
    mem_a[1731] = 8'b00000000;
    mem_a[1732] = 8'b00000000;
    mem_a[1733] = 8'b11100000;
    mem_a[1734] = 8'b11111111;
    mem_a[1735] = 8'b11111111;
    mem_a[1736] = 8'b11111111;
    mem_a[1737] = 8'b11111111;
    mem_a[1738] = 8'b11111111;
    mem_a[1739] = 8'b00000111;
    mem_a[1740] = 8'b00000000;
    mem_a[1741] = 8'b00000000;
    mem_a[1742] = 8'b00000000;
    mem_a[1743] = 8'b00000000;
    mem_a[1744] = 8'b00000000;
    mem_a[1745] = 8'b00000000;
    mem_a[1746] = 8'b00000000;
    mem_a[1747] = 8'b00000000;
    mem_a[1748] = 8'b00000000;
    mem_a[1749] = 8'b11110000;
    mem_a[1750] = 8'b11111111;
    mem_a[1751] = 8'b11111111;
    mem_a[1752] = 8'b11111111;
    mem_a[1753] = 8'b11111111;
    mem_a[1754] = 8'b11111111;
    mem_a[1755] = 8'b00000111;
    mem_a[1756] = 8'b00000000;
    mem_a[1757] = 8'b00000000;
    mem_a[1758] = 8'b00000000;
    mem_a[1759] = 8'b00000000;
    mem_a[1760] = 8'b00000000;
    mem_a[1761] = 8'b00000000;
    mem_a[1762] = 8'b00000000;
    mem_a[1763] = 8'b00000000;
    mem_a[1764] = 8'b00000000;
    mem_a[1765] = 8'b11110000;
    mem_a[1766] = 8'b11111111;
    mem_a[1767] = 8'b11111111;
    mem_a[1768] = 8'b11111111;
    mem_a[1769] = 8'b11111111;
    mem_a[1770] = 8'b11111111;
    mem_a[1771] = 8'b00000111;
    mem_a[1772] = 8'b00000000;
    mem_a[1773] = 8'b00000000;
    mem_a[1774] = 8'b00000000;
    mem_a[1775] = 8'b00000000;
    mem_a[1776] = 8'b00000000;
    mem_a[1777] = 8'b00000000;
    mem_a[1778] = 8'b00000000;
    mem_a[1779] = 8'b00000000;
    mem_a[1780] = 8'b00000000;
    mem_a[1781] = 8'b00000000;
    mem_a[1782] = 8'b11111110;
    mem_a[1783] = 8'b11111111;
    mem_a[1784] = 8'b11111111;
    mem_a[1785] = 8'b11111111;
    mem_a[1786] = 8'b11111111;
    mem_a[1787] = 8'b00001111;
    mem_a[1788] = 8'b00000000;
    mem_a[1789] = 8'b00000000;
    mem_a[1790] = 8'b00000000;
    mem_a[1791] = 8'b00000000;
    mem_a[1792] = 8'b00000000;
    mem_a[1793] = 8'b00000000;
    mem_a[1794] = 8'b00000000;
    mem_a[1795] = 8'b00000000;
    mem_a[1796] = 8'b00000000;
    mem_a[1797] = 8'b00000000;
    mem_a[1798] = 8'b11111100;
    mem_a[1799] = 8'b11111111;
    mem_a[1800] = 8'b11111111;
    mem_a[1801] = 8'b11111111;
    mem_a[1802] = 8'b11111111;
    mem_a[1803] = 8'b00001111;
    mem_a[1804] = 8'b00000000;
    mem_a[1805] = 8'b00000000;
    mem_a[1806] = 8'b00000000;
    mem_a[1807] = 8'b00000000;
    mem_a[1808] = 8'b00000000;
    mem_a[1809] = 8'b00000000;
    mem_a[1810] = 8'b00000000;
    mem_a[1811] = 8'b00000000;
    mem_a[1812] = 8'b00000000;
    mem_a[1813] = 8'b00000000;
    mem_a[1814] = 8'b11111100;
    mem_a[1815] = 8'b11111111;
    mem_a[1816] = 8'b11111111;
    mem_a[1817] = 8'b11111111;
    mem_a[1818] = 8'b11111111;
    mem_a[1819] = 8'b00001111;
    mem_a[1820] = 8'b00000000;
    mem_a[1821] = 8'b00000000;
    mem_a[1822] = 8'b00000000;
    mem_a[1823] = 8'b00000000;
    mem_a[1824] = 8'b00000000;
    mem_a[1825] = 8'b00000000;
    mem_a[1826] = 8'b00000000;
    mem_a[1827] = 8'b00000000;
    mem_a[1828] = 8'b00000000;
    mem_a[1829] = 8'b00000000;
    mem_a[1830] = 8'b11111100;
    mem_a[1831] = 8'b11111111;
    mem_a[1832] = 8'b11111111;
    mem_a[1833] = 8'b11111111;
    mem_a[1834] = 8'b11111111;
    mem_a[1835] = 8'b00011111;
    mem_a[1836] = 8'b00000000;
    mem_a[1837] = 8'b00000000;
    mem_a[1838] = 8'b00000000;
    mem_a[1839] = 8'b00000000;
    mem_a[1840] = 8'b00000000;
    mem_a[1841] = 8'b00000000;
    mem_a[1842] = 8'b00000000;
    mem_a[1843] = 8'b00000000;
    mem_a[1844] = 8'b00000000;
    mem_a[1845] = 8'b00000000;
    mem_a[1846] = 8'b11111110;
    mem_a[1847] = 8'b11111111;
    mem_a[1848] = 8'b11111111;
    mem_a[1849] = 8'b11111111;
    mem_a[1850] = 8'b11111111;
    mem_a[1851] = 8'b00011111;
    mem_a[1852] = 8'b00000000;
    mem_a[1853] = 8'b00000000;
    mem_a[1854] = 8'b00000000;
    mem_a[1855] = 8'b00000000;
    mem_a[1856] = 8'b00000000;
    mem_a[1857] = 8'b00000000;
    mem_a[1858] = 8'b00000000;
    mem_a[1859] = 8'b00000000;
    mem_a[1860] = 8'b00000000;
    mem_a[1861] = 8'b00000000;
    mem_a[1862] = 8'b11111110;
    mem_a[1863] = 8'b11111111;
    mem_a[1864] = 8'b11111111;
    mem_a[1865] = 8'b11111111;
    mem_a[1866] = 8'b11111111;
    mem_a[1867] = 8'b00011111;
    mem_a[1868] = 8'b00000000;
    mem_a[1869] = 8'b00000000;
    mem_a[1870] = 8'b00000000;
    mem_a[1871] = 8'b00000000;
    mem_a[1872] = 8'b00000000;
    mem_a[1873] = 8'b00000000;
    mem_a[1874] = 8'b00000000;
    mem_a[1875] = 8'b00000000;
    mem_a[1876] = 8'b00000000;
    mem_a[1877] = 8'b00000000;
    mem_a[1878] = 8'b11111111;
    mem_a[1879] = 8'b11111111;
    mem_a[1880] = 8'b11111111;
    mem_a[1881] = 8'b11111111;
    mem_a[1882] = 8'b11111111;
    mem_a[1883] = 8'b00111111;
    mem_a[1884] = 8'b00000000;
    mem_a[1885] = 8'b00000000;
    mem_a[1886] = 8'b00000000;
    mem_a[1887] = 8'b00000000;
    mem_a[1888] = 8'b00000000;
    mem_a[1889] = 8'b00000000;
    mem_a[1890] = 8'b00000000;
    mem_a[1891] = 8'b00000000;
    mem_a[1892] = 8'b00000000;
    mem_a[1893] = 8'b00000000;
    mem_a[1894] = 8'b11111111;
    mem_a[1895] = 8'b11111111;
    mem_a[1896] = 8'b11111111;
    mem_a[1897] = 8'b11111111;
    mem_a[1898] = 8'b11111111;
    mem_a[1899] = 8'b00111111;
    mem_a[1900] = 8'b00000000;
    mem_a[1901] = 8'b00000000;
    mem_a[1902] = 8'b00000000;
    mem_a[1903] = 8'b00000000;
    mem_a[1904] = 8'b00000000;
    mem_a[1905] = 8'b00000000;
    mem_a[1906] = 8'b00000000;
    mem_a[1907] = 8'b00000000;
    mem_a[1908] = 8'b00000000;
    mem_a[1909] = 8'b10000000;
    mem_a[1910] = 8'b11111111;
    mem_a[1911] = 8'b11111111;
    mem_a[1912] = 8'b11111111;
    mem_a[1913] = 8'b11111111;
    mem_a[1914] = 8'b11111111;
    mem_a[1915] = 8'b00111111;
    mem_a[1916] = 8'b00000000;
    mem_a[1917] = 8'b00000000;
    mem_a[1918] = 8'b00000000;
    mem_a[1919] = 8'b00000000;
    mem_a[1920] = 8'b00000000;
    mem_a[1921] = 8'b00000000;
    mem_a[1922] = 8'b00000000;
    mem_a[1923] = 8'b00000000;
    mem_a[1924] = 8'b00000000;
    mem_a[1925] = 8'b10000000;
    mem_a[1926] = 8'b11111111;
    mem_a[1927] = 8'b11111111;
    mem_a[1928] = 8'b11111111;
    mem_a[1929] = 8'b11111111;
    mem_a[1930] = 8'b11111111;
    mem_a[1931] = 8'b00111111;
    mem_a[1932] = 8'b00000000;
    mem_a[1933] = 8'b00000000;
    mem_a[1934] = 8'b00000000;
    mem_a[1935] = 8'b00000000;
    mem_a[1936] = 8'b00000000;
    mem_a[1937] = 8'b00000000;
    mem_a[1938] = 8'b00000000;
    mem_a[1939] = 8'b00000000;
    mem_a[1940] = 8'b00000000;
    mem_a[1941] = 8'b10000000;
    mem_a[1942] = 8'b11111111;
    mem_a[1943] = 8'b11111111;
    mem_a[1944] = 8'b11111111;
    mem_a[1945] = 8'b11111111;
    mem_a[1946] = 8'b11111111;
    mem_a[1947] = 8'b00111111;
    mem_a[1948] = 8'b00000000;
    mem_a[1949] = 8'b00000000;
    mem_a[1950] = 8'b00000000;
    mem_a[1951] = 8'b00000000;
    mem_a[1952] = 8'b00000000;
    mem_a[1953] = 8'b00000000;
    mem_a[1954] = 8'b00000000;
    mem_a[1955] = 8'b00000000;
    mem_a[1956] = 8'b00000000;
    mem_a[1957] = 8'b11000000;
    mem_a[1958] = 8'b11111111;
    mem_a[1959] = 8'b11111111;
    mem_a[1960] = 8'b11111111;
    mem_a[1961] = 8'b11111111;
    mem_a[1962] = 8'b11111111;
    mem_a[1963] = 8'b01111111;
    mem_a[1964] = 8'b00000000;
    mem_a[1965] = 8'b00000000;
    mem_a[1966] = 8'b00000000;
    mem_a[1967] = 8'b00000000;
    mem_a[1968] = 8'b00000000;
    mem_a[1969] = 8'b00000000;
    mem_a[1970] = 8'b00000000;
    mem_a[1971] = 8'b00000000;
    mem_a[1972] = 8'b00000000;
    mem_a[1973] = 8'b11000000;
    mem_a[1974] = 8'b11111111;
    mem_a[1975] = 8'b11111111;
    mem_a[1976] = 8'b11111111;
    mem_a[1977] = 8'b11111111;
    mem_a[1978] = 8'b11111111;
    mem_a[1979] = 8'b01111111;
    mem_a[1980] = 8'b00000000;
    mem_a[1981] = 8'b00000000;
    mem_a[1982] = 8'b00000000;
    mem_a[1983] = 8'b00000000;
    mem_a[1984] = 8'b00000000;
    mem_a[1985] = 8'b00000000;
    mem_a[1986] = 8'b00000000;
    mem_a[1987] = 8'b00000000;
    mem_a[1988] = 8'b00000000;
    mem_a[1989] = 8'b11000000;
    mem_a[1990] = 8'b11111111;
    mem_a[1991] = 8'b11111111;
    mem_a[1992] = 8'b11111111;
    mem_a[1993] = 8'b11111111;
    mem_a[1994] = 8'b11111111;
    mem_a[1995] = 8'b01111111;
    mem_a[1996] = 8'b00000000;
    mem_a[1997] = 8'b00000000;
    mem_a[1998] = 8'b00000000;
    mem_a[1999] = 8'b00000000;
    mem_a[2000] = 8'b00000000;
    mem_a[2001] = 8'b00000000;
    mem_a[2002] = 8'b00000000;
    mem_a[2003] = 8'b00000000;
    mem_a[2004] = 8'b00000000;
    mem_a[2005] = 8'b11000000;
    mem_a[2006] = 8'b11111111;
    mem_a[2007] = 8'b11111111;
    mem_a[2008] = 8'b11111111;
    mem_a[2009] = 8'b11111111;
    mem_a[2010] = 8'b11111111;
    mem_a[2011] = 8'b01111111;
    mem_a[2012] = 8'b00000000;
    mem_a[2013] = 8'b00000000;
    mem_a[2014] = 8'b00000000;
    mem_a[2015] = 8'b00000000;
    mem_a[2016] = 8'b00000000;
    mem_a[2017] = 8'b00000000;
    mem_a[2018] = 8'b00000000;
    mem_a[2019] = 8'b00000000;
    mem_a[2020] = 8'b00000000;
    mem_a[2021] = 8'b11000000;
    mem_a[2022] = 8'b11111111;
    mem_a[2023] = 8'b11111111;
    mem_a[2024] = 8'b11111111;
    mem_a[2025] = 8'b11111111;
    mem_a[2026] = 8'b11111111;
    mem_a[2027] = 8'b01111111;
    mem_a[2028] = 8'b00000000;
    mem_a[2029] = 8'b00000000;
    mem_a[2030] = 8'b00000000;
    mem_a[2031] = 8'b00000000;
    mem_a[2032] = 8'b00000000;
    mem_a[2033] = 8'b00000000;
    mem_a[2034] = 8'b00000000;
    mem_a[2035] = 8'b00000000;
    mem_a[2036] = 8'b00000000;
    mem_a[2037] = 8'b11111000;
    mem_a[2038] = 8'b11111111;
    mem_a[2039] = 8'b11111111;
    mem_a[2040] = 8'b11111111;
    mem_a[2041] = 8'b11111111;
    mem_a[2042] = 8'b11111111;
    mem_a[2043] = 8'b11111111;
    mem_a[2044] = 8'b00000011;
    mem_a[2045] = 8'b00000000;
    mem_a[2046] = 8'b00000000;
    mem_a[2047] = 8'b00000000;
end

reg [7:0] mem_b [0:2047];
initial begin
    mem_b[0] = 8'b00000000;
    mem_b[1] = 8'b00000000;
    mem_b[2] = 8'b00000000;
    mem_b[3] = 8'b00000000;
    mem_b[4] = 8'b00000000;
    mem_b[5] = 8'b00000000;
    mem_b[6] = 8'b00000000;
    mem_b[7] = 8'b00000000;
    mem_b[8] = 8'b00000000;
    mem_b[9] = 8'b00000000;
    mem_b[10] = 8'b00000000;
    mem_b[11] = 8'b00000000;
    mem_b[12] = 8'b00000000;
    mem_b[13] = 8'b00000000;
    mem_b[14] = 8'b00000000;
    mem_b[15] = 8'b00000000;
    mem_b[16] = 8'b00000000;
    mem_b[17] = 8'b00000000;
    mem_b[18] = 8'b00000000;
    mem_b[19] = 8'b00000000;
    mem_b[20] = 8'b00000000;
    mem_b[21] = 8'b00000000;
    mem_b[22] = 8'b00000000;
    mem_b[23] = 8'b00000000;
    mem_b[24] = 8'b00000000;
    mem_b[25] = 8'b00000000;
    mem_b[26] = 8'b00000000;
    mem_b[27] = 8'b00000000;
    mem_b[28] = 8'b00000000;
    mem_b[29] = 8'b11111000;
    mem_b[30] = 8'b00000000;
    mem_b[31] = 8'b00000000;
    mem_b[32] = 8'b00000000;
    mem_b[33] = 8'b10000000;
    mem_b[34] = 8'b00001111;
    mem_b[35] = 8'b00000000;
    mem_b[36] = 8'b00000000;
    mem_b[37] = 8'b00000000;
    mem_b[38] = 8'b00000000;
    mem_b[39] = 8'b00000000;
    mem_b[40] = 8'b00000000;
    mem_b[41] = 8'b00000000;
    mem_b[42] = 8'b00000000;
    mem_b[43] = 8'b00000000;
    mem_b[44] = 8'b00000000;
    mem_b[45] = 8'b11111111;
    mem_b[46] = 8'b00000000;
    mem_b[47] = 8'b00000000;
    mem_b[48] = 8'b00000000;
    mem_b[49] = 8'b10000000;
    mem_b[50] = 8'b11111111;
    mem_b[51] = 8'b00000000;
    mem_b[52] = 8'b00000000;
    mem_b[53] = 8'b00000000;
    mem_b[54] = 8'b00000000;
    mem_b[55] = 8'b00000000;
    mem_b[56] = 8'b00000000;
    mem_b[57] = 8'b00000000;
    mem_b[58] = 8'b00000000;
    mem_b[59] = 8'b00000000;
    mem_b[60] = 8'b11000000;
    mem_b[61] = 8'b11111111;
    mem_b[62] = 8'b00000001;
    mem_b[63] = 8'b00000000;
    mem_b[64] = 8'b00000000;
    mem_b[65] = 8'b10000000;
    mem_b[66] = 8'b11111111;
    mem_b[67] = 8'b00000111;
    mem_b[68] = 8'b00000000;
    mem_b[69] = 8'b00000000;
    mem_b[70] = 8'b00000000;
    mem_b[71] = 8'b00000000;
    mem_b[72] = 8'b00000000;
    mem_b[73] = 8'b00000000;
    mem_b[74] = 8'b00000000;
    mem_b[75] = 8'b00000000;
    mem_b[76] = 8'b11111000;
    mem_b[77] = 8'b11111111;
    mem_b[78] = 8'b00000001;
    mem_b[79] = 8'b00000000;
    mem_b[80] = 8'b00000000;
    mem_b[81] = 8'b10000000;
    mem_b[82] = 8'b11111111;
    mem_b[83] = 8'b00011111;
    mem_b[84] = 8'b00000000;
    mem_b[85] = 8'b00000000;
    mem_b[86] = 8'b00000000;
    mem_b[87] = 8'b00000000;
    mem_b[88] = 8'b00000000;
    mem_b[89] = 8'b00000000;
    mem_b[90] = 8'b00000000;
    mem_b[91] = 8'b00000000;
    mem_b[92] = 8'b11111110;
    mem_b[93] = 8'b11111111;
    mem_b[94] = 8'b00000001;
    mem_b[95] = 8'b00000000;
    mem_b[96] = 8'b00000000;
    mem_b[97] = 8'b11000000;
    mem_b[98] = 8'b11111111;
    mem_b[99] = 8'b00111111;
    mem_b[100] = 8'b00000000;
    mem_b[101] = 8'b00000000;
    mem_b[102] = 8'b00000000;
    mem_b[103] = 8'b00000000;
    mem_b[104] = 8'b00000000;
    mem_b[105] = 8'b00000000;
    mem_b[106] = 8'b00000000;
    mem_b[107] = 8'b10000000;
    mem_b[108] = 8'b11111111;
    mem_b[109] = 8'b11111111;
    mem_b[110] = 8'b00000011;
    mem_b[111] = 8'b00000000;
    mem_b[112] = 8'b00000000;
    mem_b[113] = 8'b11000000;
    mem_b[114] = 8'b11111111;
    mem_b[115] = 8'b01111111;
    mem_b[116] = 8'b00000000;
    mem_b[117] = 8'b00000000;
    mem_b[118] = 8'b00000000;
    mem_b[119] = 8'b00000000;
    mem_b[120] = 8'b00000000;
    mem_b[121] = 8'b00000000;
    mem_b[122] = 8'b00000000;
    mem_b[123] = 8'b11100000;
    mem_b[124] = 8'b11111111;
    mem_b[125] = 8'b11111111;
    mem_b[126] = 8'b00000011;
    mem_b[127] = 8'b00000000;
    mem_b[128] = 8'b00000000;
    mem_b[129] = 8'b11000000;
    mem_b[130] = 8'b11111111;
    mem_b[131] = 8'b11111111;
    mem_b[132] = 8'b00000000;
    mem_b[133] = 8'b00000000;
    mem_b[134] = 8'b00000000;
    mem_b[135] = 8'b00000000;
    mem_b[136] = 8'b00000000;
    mem_b[137] = 8'b00000000;
    mem_b[138] = 8'b00000000;
    mem_b[139] = 8'b11110000;
    mem_b[140] = 8'b11111111;
    mem_b[141] = 8'b11111111;
    mem_b[142] = 8'b00000011;
    mem_b[143] = 8'b00000000;
    mem_b[144] = 8'b00000000;
    mem_b[145] = 8'b11000000;
    mem_b[146] = 8'b11111111;
    mem_b[147] = 8'b11111111;
    mem_b[148] = 8'b00000001;
    mem_b[149] = 8'b00000000;
    mem_b[150] = 8'b00001110;
    mem_b[151] = 8'b00000000;
    mem_b[152] = 8'b00000000;
    mem_b[153] = 8'b00000000;
    mem_b[154] = 8'b00000000;
    mem_b[155] = 8'b11111100;
    mem_b[156] = 8'b11111111;
    mem_b[157] = 8'b11111111;
    mem_b[158] = 8'b00000111;
    mem_b[159] = 8'b00000000;
    mem_b[160] = 8'b00000000;
    mem_b[161] = 8'b11100000;
    mem_b[162] = 8'b11111111;
    mem_b[163] = 8'b11111111;
    mem_b[164] = 8'b00000111;
    mem_b[165] = 8'b00000000;
    mem_b[166] = 8'b11111110;
    mem_b[167] = 8'b00001111;
    mem_b[168] = 8'b00000000;
    mem_b[169] = 8'b00000000;
    mem_b[170] = 8'b00000000;
    mem_b[171] = 8'b11111110;
    mem_b[172] = 8'b11111111;
    mem_b[173] = 8'b11111111;
    mem_b[174] = 8'b00000111;
    mem_b[175] = 8'b00000000;
    mem_b[176] = 8'b00000000;
    mem_b[177] = 8'b11100000;
    mem_b[178] = 8'b11111111;
    mem_b[179] = 8'b11111111;
    mem_b[180] = 8'b00001111;
    mem_b[181] = 8'b00000000;
    mem_b[182] = 8'b11111110;
    mem_b[183] = 8'b01111111;
    mem_b[184] = 8'b00000000;
    mem_b[185] = 8'b00000000;
    mem_b[186] = 8'b00000000;
    mem_b[187] = 8'b11111111;
    mem_b[188] = 8'b11111111;
    mem_b[189] = 8'b11111111;
    mem_b[190] = 8'b00000111;
    mem_b[191] = 8'b00000000;
    mem_b[192] = 8'b00000000;
    mem_b[193] = 8'b11100000;
    mem_b[194] = 8'b11111111;
    mem_b[195] = 8'b11111111;
    mem_b[196] = 8'b00111111;
    mem_b[197] = 8'b00000000;
    mem_b[198] = 8'b11111110;
    mem_b[199] = 8'b11111111;
    mem_b[200] = 8'b00000011;
    mem_b[201] = 8'b00000000;
    mem_b[202] = 8'b11000000;
    mem_b[203] = 8'b11111111;
    mem_b[204] = 8'b11111111;
    mem_b[205] = 8'b11111111;
    mem_b[206] = 8'b00001111;
    mem_b[207] = 8'b00000000;
    mem_b[208] = 8'b00000000;
    mem_b[209] = 8'b11100000;
    mem_b[210] = 8'b11111111;
    mem_b[211] = 8'b11111111;
    mem_b[212] = 8'b01111111;
    mem_b[213] = 8'b00000000;
    mem_b[214] = 8'b11111110;
    mem_b[215] = 8'b11111111;
    mem_b[216] = 8'b00011111;
    mem_b[217] = 8'b00000000;
    mem_b[218] = 8'b11100000;
    mem_b[219] = 8'b11111111;
    mem_b[220] = 8'b11111111;
    mem_b[221] = 8'b11111111;
    mem_b[222] = 8'b00001111;
    mem_b[223] = 8'b00000000;
    mem_b[224] = 8'b00000000;
    mem_b[225] = 8'b11100000;
    mem_b[226] = 8'b11111111;
    mem_b[227] = 8'b11111111;
    mem_b[228] = 8'b11111111;
    mem_b[229] = 8'b00000000;
    mem_b[230] = 8'b11111100;
    mem_b[231] = 8'b11111111;
    mem_b[232] = 8'b01111111;
    mem_b[233] = 8'b00000000;
    mem_b[234] = 8'b11100000;
    mem_b[235] = 8'b11111111;
    mem_b[236] = 8'b11111111;
    mem_b[237] = 8'b11111111;
    mem_b[238] = 8'b00001111;
    mem_b[239] = 8'b00000000;
    mem_b[240] = 8'b00000000;
    mem_b[241] = 8'b11110000;
    mem_b[242] = 8'b11111111;
    mem_b[243] = 8'b11111111;
    mem_b[244] = 8'b11111111;
    mem_b[245] = 8'b00000001;
    mem_b[246] = 8'b11111100;
    mem_b[247] = 8'b11111111;
    mem_b[248] = 8'b11111111;
    mem_b[249] = 8'b00000001;
    mem_b[250] = 8'b11110000;
    mem_b[251] = 8'b11111111;
    mem_b[252] = 8'b11111111;
    mem_b[253] = 8'b11111111;
    mem_b[254] = 8'b00001111;
    mem_b[255] = 8'b00000000;
    mem_b[256] = 8'b00000000;
    mem_b[257] = 8'b11110000;
    mem_b[258] = 8'b11111111;
    mem_b[259] = 8'b11111111;
    mem_b[260] = 8'b11111111;
    mem_b[261] = 8'b00000011;
    mem_b[262] = 8'b11111100;
    mem_b[263] = 8'b11111111;
    mem_b[264] = 8'b11111111;
    mem_b[265] = 8'b00000111;
    mem_b[266] = 8'b11110000;
    mem_b[267] = 8'b11111111;
    mem_b[268] = 8'b11111111;
    mem_b[269] = 8'b11111111;
    mem_b[270] = 8'b00011111;
    mem_b[271] = 8'b00000000;
    mem_b[272] = 8'b00000000;
    mem_b[273] = 8'b11110000;
    mem_b[274] = 8'b11111111;
    mem_b[275] = 8'b11111111;
    mem_b[276] = 8'b11111111;
    mem_b[277] = 8'b00000111;
    mem_b[278] = 8'b11111000;
    mem_b[279] = 8'b11111111;
    mem_b[280] = 8'b11111111;
    mem_b[281] = 8'b00001111;
    mem_b[282] = 8'b11111000;
    mem_b[283] = 8'b11111111;
    mem_b[284] = 8'b11111111;
    mem_b[285] = 8'b11111111;
    mem_b[286] = 8'b00011111;
    mem_b[287] = 8'b00000000;
    mem_b[288] = 8'b00000000;
    mem_b[289] = 8'b11110000;
    mem_b[290] = 8'b11111111;
    mem_b[291] = 8'b11111111;
    mem_b[292] = 8'b11111111;
    mem_b[293] = 8'b00000111;
    mem_b[294] = 8'b11111000;
    mem_b[295] = 8'b11111111;
    mem_b[296] = 8'b11111111;
    mem_b[297] = 8'b00011111;
    mem_b[298] = 8'b11111100;
    mem_b[299] = 8'b11111111;
    mem_b[300] = 8'b11111111;
    mem_b[301] = 8'b11111111;
    mem_b[302] = 8'b00011111;
    mem_b[303] = 8'b00000000;
    mem_b[304] = 8'b00000000;
    mem_b[305] = 8'b11110000;
    mem_b[306] = 8'b11111111;
    mem_b[307] = 8'b11111111;
    mem_b[308] = 8'b11111111;
    mem_b[309] = 8'b00001111;
    mem_b[310] = 8'b11111000;
    mem_b[311] = 8'b11111111;
    mem_b[312] = 8'b11111111;
    mem_b[313] = 8'b00111111;
    mem_b[314] = 8'b11111100;
    mem_b[315] = 8'b11111111;
    mem_b[316] = 8'b11111111;
    mem_b[317] = 8'b11111111;
    mem_b[318] = 8'b00011111;
    mem_b[319] = 8'b00000000;
    mem_b[320] = 8'b00000000;
    mem_b[321] = 8'b11111000;
    mem_b[322] = 8'b11111111;
    mem_b[323] = 8'b11111111;
    mem_b[324] = 8'b11111111;
    mem_b[325] = 8'b00011111;
    mem_b[326] = 8'b11110000;
    mem_b[327] = 8'b11111111;
    mem_b[328] = 8'b11111111;
    mem_b[329] = 8'b11111111;
    mem_b[330] = 8'b11111110;
    mem_b[331] = 8'b11111111;
    mem_b[332] = 8'b11111111;
    mem_b[333] = 8'b11111111;
    mem_b[334] = 8'b00011111;
    mem_b[335] = 8'b00000000;
    mem_b[336] = 8'b00000000;
    mem_b[337] = 8'b11111000;
    mem_b[338] = 8'b11111111;
    mem_b[339] = 8'b11111111;
    mem_b[340] = 8'b11111111;
    mem_b[341] = 8'b00111111;
    mem_b[342] = 8'b11110000;
    mem_b[343] = 8'b11111111;
    mem_b[344] = 8'b11111111;
    mem_b[345] = 8'b11111111;
    mem_b[346] = 8'b11111111;
    mem_b[347] = 8'b11111111;
    mem_b[348] = 8'b11111111;
    mem_b[349] = 8'b11111111;
    mem_b[350] = 8'b00111111;
    mem_b[351] = 8'b00000000;
    mem_b[352] = 8'b00000000;
    mem_b[353] = 8'b11111000;
    mem_b[354] = 8'b11111111;
    mem_b[355] = 8'b11111111;
    mem_b[356] = 8'b11111111;
    mem_b[357] = 8'b01111111;
    mem_b[358] = 8'b11100000;
    mem_b[359] = 8'b11111111;
    mem_b[360] = 8'b11111111;
    mem_b[361] = 8'b11111111;
    mem_b[362] = 8'b11111111;
    mem_b[363] = 8'b11111111;
    mem_b[364] = 8'b11111111;
    mem_b[365] = 8'b11111111;
    mem_b[366] = 8'b00111111;
    mem_b[367] = 8'b00000000;
    mem_b[368] = 8'b00000000;
    mem_b[369] = 8'b11111000;
    mem_b[370] = 8'b11111111;
    mem_b[371] = 8'b11111111;
    mem_b[372] = 8'b11111111;
    mem_b[373] = 8'b11111111;
    mem_b[374] = 8'b11000000;
    mem_b[375] = 8'b11111111;
    mem_b[376] = 8'b11111111;
    mem_b[377] = 8'b11111111;
    mem_b[378] = 8'b11111111;
    mem_b[379] = 8'b11111111;
    mem_b[380] = 8'b11111111;
    mem_b[381] = 8'b11111111;
    mem_b[382] = 8'b00111111;
    mem_b[383] = 8'b00000000;
    mem_b[384] = 8'b00000000;
    mem_b[385] = 8'b11111000;
    mem_b[386] = 8'b11111111;
    mem_b[387] = 8'b11111111;
    mem_b[388] = 8'b11111111;
    mem_b[389] = 8'b11111111;
    mem_b[390] = 8'b10000001;
    mem_b[391] = 8'b11111111;
    mem_b[392] = 8'b11111111;
    mem_b[393] = 8'b11111111;
    mem_b[394] = 8'b11111111;
    mem_b[395] = 8'b11111111;
    mem_b[396] = 8'b11111111;
    mem_b[397] = 8'b11111111;
    mem_b[398] = 8'b00111111;
    mem_b[399] = 8'b00000000;
    mem_b[400] = 8'b00000000;
    mem_b[401] = 8'b11111000;
    mem_b[402] = 8'b11111111;
    mem_b[403] = 8'b11111111;
    mem_b[404] = 8'b11111111;
    mem_b[405] = 8'b11111111;
    mem_b[406] = 8'b11110011;
    mem_b[407] = 8'b11111111;
    mem_b[408] = 8'b11111111;
    mem_b[409] = 8'b11111111;
    mem_b[410] = 8'b11111111;
    mem_b[411] = 8'b11111111;
    mem_b[412] = 8'b11111111;
    mem_b[413] = 8'b11111111;
    mem_b[414] = 8'b01111111;
    mem_b[415] = 8'b00000000;
    mem_b[416] = 8'b00000000;
    mem_b[417] = 8'b11111000;
    mem_b[418] = 8'b11111111;
    mem_b[419] = 8'b11111111;
    mem_b[420] = 8'b11111111;
    mem_b[421] = 8'b11111111;
    mem_b[422] = 8'b11111111;
    mem_b[423] = 8'b11111111;
    mem_b[424] = 8'b11111111;
    mem_b[425] = 8'b11111111;
    mem_b[426] = 8'b11111111;
    mem_b[427] = 8'b11111111;
    mem_b[428] = 8'b11111111;
    mem_b[429] = 8'b11111111;
    mem_b[430] = 8'b01111111;
    mem_b[431] = 8'b00000000;
    mem_b[432] = 8'b00000000;
    mem_b[433] = 8'b11111000;
    mem_b[434] = 8'b11111111;
    mem_b[435] = 8'b11111111;
    mem_b[436] = 8'b11111111;
    mem_b[437] = 8'b11111111;
    mem_b[438] = 8'b11111111;
    mem_b[439] = 8'b11111111;
    mem_b[440] = 8'b11111111;
    mem_b[441] = 8'b11111111;
    mem_b[442] = 8'b11111111;
    mem_b[443] = 8'b11111111;
    mem_b[444] = 8'b11111111;
    mem_b[445] = 8'b11111111;
    mem_b[446] = 8'b01111111;
    mem_b[447] = 8'b00000000;
    mem_b[448] = 8'b00000000;
    mem_b[449] = 8'b11111100;
    mem_b[450] = 8'b11111111;
    mem_b[451] = 8'b11111111;
    mem_b[452] = 8'b11111111;
    mem_b[453] = 8'b11111111;
    mem_b[454] = 8'b11111111;
    mem_b[455] = 8'b11111111;
    mem_b[456] = 8'b11111111;
    mem_b[457] = 8'b11111111;
    mem_b[458] = 8'b11111111;
    mem_b[459] = 8'b11111111;
    mem_b[460] = 8'b11111111;
    mem_b[461] = 8'b11111111;
    mem_b[462] = 8'b01111111;
    mem_b[463] = 8'b00000000;
    mem_b[464] = 8'b00000000;
    mem_b[465] = 8'b11111100;
    mem_b[466] = 8'b11111111;
    mem_b[467] = 8'b11111111;
    mem_b[468] = 8'b11111111;
    mem_b[469] = 8'b11111111;
    mem_b[470] = 8'b11111111;
    mem_b[471] = 8'b11111111;
    mem_b[472] = 8'b11111111;
    mem_b[473] = 8'b11111111;
    mem_b[474] = 8'b11111111;
    mem_b[475] = 8'b11111111;
    mem_b[476] = 8'b11111111;
    mem_b[477] = 8'b11111111;
    mem_b[478] = 8'b01111111;
    mem_b[479] = 8'b00000000;
    mem_b[480] = 8'b00000000;
    mem_b[481] = 8'b11111100;
    mem_b[482] = 8'b11111111;
    mem_b[483] = 8'b11111111;
    mem_b[484] = 8'b11111111;
    mem_b[485] = 8'b11111111;
    mem_b[486] = 8'b11111111;
    mem_b[487] = 8'b11111111;
    mem_b[488] = 8'b11111111;
    mem_b[489] = 8'b11111111;
    mem_b[490] = 8'b11111111;
    mem_b[491] = 8'b11111111;
    mem_b[492] = 8'b11111111;
    mem_b[493] = 8'b11111111;
    mem_b[494] = 8'b01111111;
    mem_b[495] = 8'b00000000;
    mem_b[496] = 8'b00000000;
    mem_b[497] = 8'b11111100;
    mem_b[498] = 8'b11111111;
    mem_b[499] = 8'b11111111;
    mem_b[500] = 8'b11111111;
    mem_b[501] = 8'b11111111;
    mem_b[502] = 8'b11111111;
    mem_b[503] = 8'b11111111;
    mem_b[504] = 8'b11111111;
    mem_b[505] = 8'b11111111;
    mem_b[506] = 8'b11111111;
    mem_b[507] = 8'b11111111;
    mem_b[508] = 8'b11111111;
    mem_b[509] = 8'b11111111;
    mem_b[510] = 8'b11111111;
    mem_b[511] = 8'b00000000;
    mem_b[512] = 8'b00000000;
    mem_b[513] = 8'b11111100;
    mem_b[514] = 8'b11111111;
    mem_b[515] = 8'b11111111;
    mem_b[516] = 8'b11111111;
    mem_b[517] = 8'b11111111;
    mem_b[518] = 8'b11111111;
    mem_b[519] = 8'b11111111;
    mem_b[520] = 8'b11111111;
    mem_b[521] = 8'b11111111;
    mem_b[522] = 8'b11111111;
    mem_b[523] = 8'b11111111;
    mem_b[524] = 8'b11111111;
    mem_b[525] = 8'b11111111;
    mem_b[526] = 8'b11111111;
    mem_b[527] = 8'b00000000;
    mem_b[528] = 8'b00000000;
    mem_b[529] = 8'b11111100;
    mem_b[530] = 8'b11111111;
    mem_b[531] = 8'b11111111;
    mem_b[532] = 8'b11111111;
    mem_b[533] = 8'b11111111;
    mem_b[534] = 8'b11111111;
    mem_b[535] = 8'b11111111;
    mem_b[536] = 8'b11111111;
    mem_b[537] = 8'b11111111;
    mem_b[538] = 8'b11111111;
    mem_b[539] = 8'b11111111;
    mem_b[540] = 8'b11111111;
    mem_b[541] = 8'b11111111;
    mem_b[542] = 8'b11111111;
    mem_b[543] = 8'b00000000;
    mem_b[544] = 8'b00000000;
    mem_b[545] = 8'b11111110;
    mem_b[546] = 8'b11111111;
    mem_b[547] = 8'b11111111;
    mem_b[548] = 8'b11111111;
    mem_b[549] = 8'b11111111;
    mem_b[550] = 8'b11111111;
    mem_b[551] = 8'b11111111;
    mem_b[552] = 8'b11111111;
    mem_b[553] = 8'b11111111;
    mem_b[554] = 8'b11111111;
    mem_b[555] = 8'b11111111;
    mem_b[556] = 8'b11111111;
    mem_b[557] = 8'b11111111;
    mem_b[558] = 8'b11111111;
    mem_b[559] = 8'b00000001;
    mem_b[560] = 8'b00000000;
    mem_b[561] = 8'b11111110;
    mem_b[562] = 8'b11111111;
    mem_b[563] = 8'b11111111;
    mem_b[564] = 8'b11111111;
    mem_b[565] = 8'b11111111;
    mem_b[566] = 8'b11111111;
    mem_b[567] = 8'b11111111;
    mem_b[568] = 8'b11111111;
    mem_b[569] = 8'b11111111;
    mem_b[570] = 8'b11111111;
    mem_b[571] = 8'b11111111;
    mem_b[572] = 8'b11111111;
    mem_b[573] = 8'b11111111;
    mem_b[574] = 8'b11111111;
    mem_b[575] = 8'b00000001;
    mem_b[576] = 8'b00000000;
    mem_b[577] = 8'b11111110;
    mem_b[578] = 8'b11111111;
    mem_b[579] = 8'b11111111;
    mem_b[580] = 8'b11111111;
    mem_b[581] = 8'b11111111;
    mem_b[582] = 8'b11111111;
    mem_b[583] = 8'b11111111;
    mem_b[584] = 8'b11111111;
    mem_b[585] = 8'b11111111;
    mem_b[586] = 8'b11111111;
    mem_b[587] = 8'b11111111;
    mem_b[588] = 8'b11111111;
    mem_b[589] = 8'b11111111;
    mem_b[590] = 8'b11111111;
    mem_b[591] = 8'b00000001;
    mem_b[592] = 8'b00000000;
    mem_b[593] = 8'b11111110;
    mem_b[594] = 8'b11111111;
    mem_b[595] = 8'b11111111;
    mem_b[596] = 8'b11111111;
    mem_b[597] = 8'b11111111;
    mem_b[598] = 8'b11111111;
    mem_b[599] = 8'b11111111;
    mem_b[600] = 8'b11111111;
    mem_b[601] = 8'b11111111;
    mem_b[602] = 8'b11111111;
    mem_b[603] = 8'b11111111;
    mem_b[604] = 8'b11111111;
    mem_b[605] = 8'b11111111;
    mem_b[606] = 8'b11111111;
    mem_b[607] = 8'b00000000;
    mem_b[608] = 8'b00000000;
    mem_b[609] = 8'b11111110;
    mem_b[610] = 8'b11111111;
    mem_b[611] = 8'b11111111;
    mem_b[612] = 8'b11111111;
    mem_b[613] = 8'b11111111;
    mem_b[614] = 8'b11111111;
    mem_b[615] = 8'b11111111;
    mem_b[616] = 8'b11111111;
    mem_b[617] = 8'b11111111;
    mem_b[618] = 8'b11111111;
    mem_b[619] = 8'b11111111;
    mem_b[620] = 8'b11111111;
    mem_b[621] = 8'b11111111;
    mem_b[622] = 8'b11111111;
    mem_b[623] = 8'b00000000;
    mem_b[624] = 8'b00000000;
    mem_b[625] = 8'b11111110;
    mem_b[626] = 8'b11111111;
    mem_b[627] = 8'b11111111;
    mem_b[628] = 8'b11111111;
    mem_b[629] = 8'b11111111;
    mem_b[630] = 8'b11111111;
    mem_b[631] = 8'b11111111;
    mem_b[632] = 8'b11111111;
    mem_b[633] = 8'b11111111;
    mem_b[634] = 8'b11111111;
    mem_b[635] = 8'b11111111;
    mem_b[636] = 8'b11111111;
    mem_b[637] = 8'b11111111;
    mem_b[638] = 8'b11111111;
    mem_b[639] = 8'b00000000;
    mem_b[640] = 8'b00000000;
    mem_b[641] = 8'b11111110;
    mem_b[642] = 8'b11111111;
    mem_b[643] = 8'b11111111;
    mem_b[644] = 8'b11111111;
    mem_b[645] = 8'b11111111;
    mem_b[646] = 8'b11111111;
    mem_b[647] = 8'b11111111;
    mem_b[648] = 8'b11111111;
    mem_b[649] = 8'b11111111;
    mem_b[650] = 8'b11111111;
    mem_b[651] = 8'b11111111;
    mem_b[652] = 8'b11111111;
    mem_b[653] = 8'b11111111;
    mem_b[654] = 8'b11111111;
    mem_b[655] = 8'b00000000;
    mem_b[656] = 8'b00000000;
    mem_b[657] = 8'b11111110;
    mem_b[658] = 8'b11111111;
    mem_b[659] = 8'b11111111;
    mem_b[660] = 8'b11111111;
    mem_b[661] = 8'b11111111;
    mem_b[662] = 8'b11111111;
    mem_b[663] = 8'b11111111;
    mem_b[664] = 8'b11111111;
    mem_b[665] = 8'b11111111;
    mem_b[666] = 8'b11111111;
    mem_b[667] = 8'b11111111;
    mem_b[668] = 8'b11111111;
    mem_b[669] = 8'b11111111;
    mem_b[670] = 8'b11111111;
    mem_b[671] = 8'b00000000;
    mem_b[672] = 8'b00000000;
    mem_b[673] = 8'b11111110;
    mem_b[674] = 8'b11111111;
    mem_b[675] = 8'b11111111;
    mem_b[676] = 8'b11111111;
    mem_b[677] = 8'b11111111;
    mem_b[678] = 8'b11111111;
    mem_b[679] = 8'b11111111;
    mem_b[680] = 8'b11111111;
    mem_b[681] = 8'b11111111;
    mem_b[682] = 8'b11111111;
    mem_b[683] = 8'b11111111;
    mem_b[684] = 8'b11111111;
    mem_b[685] = 8'b11111111;
    mem_b[686] = 8'b11111111;
    mem_b[687] = 8'b00000000;
    mem_b[688] = 8'b00000000;
    mem_b[689] = 8'b11111100;
    mem_b[690] = 8'b11111111;
    mem_b[691] = 8'b11111111;
    mem_b[692] = 8'b11111111;
    mem_b[693] = 8'b11111111;
    mem_b[694] = 8'b11111111;
    mem_b[695] = 8'b11111111;
    mem_b[696] = 8'b11111111;
    mem_b[697] = 8'b11111111;
    mem_b[698] = 8'b11111111;
    mem_b[699] = 8'b11111111;
    mem_b[700] = 8'b11111111;
    mem_b[701] = 8'b11111111;
    mem_b[702] = 8'b11111111;
    mem_b[703] = 8'b00000000;
    mem_b[704] = 8'b00000000;
    mem_b[705] = 8'b11111100;
    mem_b[706] = 8'b11111111;
    mem_b[707] = 8'b11111111;
    mem_b[708] = 8'b11111111;
    mem_b[709] = 8'b11111111;
    mem_b[710] = 8'b11111111;
    mem_b[711] = 8'b11111111;
    mem_b[712] = 8'b11111111;
    mem_b[713] = 8'b11111111;
    mem_b[714] = 8'b11111111;
    mem_b[715] = 8'b11111111;
    mem_b[716] = 8'b11111111;
    mem_b[717] = 8'b11111111;
    mem_b[718] = 8'b01111111;
    mem_b[719] = 8'b00000000;
    mem_b[720] = 8'b00000000;
    mem_b[721] = 8'b11111100;
    mem_b[722] = 8'b11111111;
    mem_b[723] = 8'b11111111;
    mem_b[724] = 8'b11111111;
    mem_b[725] = 8'b11111111;
    mem_b[726] = 8'b11111111;
    mem_b[727] = 8'b11111111;
    mem_b[728] = 8'b11111111;
    mem_b[729] = 8'b11111111;
    mem_b[730] = 8'b11111111;
    mem_b[731] = 8'b11111111;
    mem_b[732] = 8'b11111111;
    mem_b[733] = 8'b11111111;
    mem_b[734] = 8'b01111111;
    mem_b[735] = 8'b00000000;
    mem_b[736] = 8'b00000000;
    mem_b[737] = 8'b11111100;
    mem_b[738] = 8'b11111111;
    mem_b[739] = 8'b11111111;
    mem_b[740] = 8'b11111111;
    mem_b[741] = 8'b11111111;
    mem_b[742] = 8'b11111111;
    mem_b[743] = 8'b11111111;
    mem_b[744] = 8'b11111111;
    mem_b[745] = 8'b11111111;
    mem_b[746] = 8'b11111111;
    mem_b[747] = 8'b11111111;
    mem_b[748] = 8'b11111111;
    mem_b[749] = 8'b11111111;
    mem_b[750] = 8'b01111111;
    mem_b[751] = 8'b00000000;
    mem_b[752] = 8'b00000000;
    mem_b[753] = 8'b11111000;
    mem_b[754] = 8'b11111111;
    mem_b[755] = 8'b11111111;
    mem_b[756] = 8'b11111111;
    mem_b[757] = 8'b11111111;
    mem_b[758] = 8'b11111111;
    mem_b[759] = 8'b11111111;
    mem_b[760] = 8'b11111111;
    mem_b[761] = 8'b11111111;
    mem_b[762] = 8'b11111111;
    mem_b[763] = 8'b11111111;
    mem_b[764] = 8'b11111111;
    mem_b[765] = 8'b11111111;
    mem_b[766] = 8'b01111111;
    mem_b[767] = 8'b00000000;
    mem_b[768] = 8'b00000000;
    mem_b[769] = 8'b11111000;
    mem_b[770] = 8'b11111111;
    mem_b[771] = 8'b11111111;
    mem_b[772] = 8'b11111111;
    mem_b[773] = 8'b11111111;
    mem_b[774] = 8'b11111111;
    mem_b[775] = 8'b11111111;
    mem_b[776] = 8'b11111111;
    mem_b[777] = 8'b11111111;
    mem_b[778] = 8'b11111111;
    mem_b[779] = 8'b11111111;
    mem_b[780] = 8'b11111111;
    mem_b[781] = 8'b11111111;
    mem_b[782] = 8'b00111111;
    mem_b[783] = 8'b00000000;
    mem_b[784] = 8'b00000000;
    mem_b[785] = 8'b11111000;
    mem_b[786] = 8'b11111111;
    mem_b[787] = 8'b11111111;
    mem_b[788] = 8'b11111111;
    mem_b[789] = 8'b11111111;
    mem_b[790] = 8'b11111111;
    mem_b[791] = 8'b11111111;
    mem_b[792] = 8'b11111111;
    mem_b[793] = 8'b11111111;
    mem_b[794] = 8'b11111111;
    mem_b[795] = 8'b11111111;
    mem_b[796] = 8'b11111111;
    mem_b[797] = 8'b11111111;
    mem_b[798] = 8'b00111111;
    mem_b[799] = 8'b00000000;
    mem_b[800] = 8'b00000000;
    mem_b[801] = 8'b11110000;
    mem_b[802] = 8'b11111111;
    mem_b[803] = 8'b11111111;
    mem_b[804] = 8'b11111111;
    mem_b[805] = 8'b11111111;
    mem_b[806] = 8'b11111111;
    mem_b[807] = 8'b11111111;
    mem_b[808] = 8'b11111111;
    mem_b[809] = 8'b11111111;
    mem_b[810] = 8'b11111111;
    mem_b[811] = 8'b11111111;
    mem_b[812] = 8'b11111111;
    mem_b[813] = 8'b11111111;
    mem_b[814] = 8'b00011111;
    mem_b[815] = 8'b00000000;
    mem_b[816] = 8'b00000000;
    mem_b[817] = 8'b11110000;
    mem_b[818] = 8'b11111111;
    mem_b[819] = 8'b11111111;
    mem_b[820] = 8'b11111111;
    mem_b[821] = 8'b11111111;
    mem_b[822] = 8'b11111111;
    mem_b[823] = 8'b11111111;
    mem_b[824] = 8'b11111111;
    mem_b[825] = 8'b11111111;
    mem_b[826] = 8'b11111111;
    mem_b[827] = 8'b11111111;
    mem_b[828] = 8'b11111111;
    mem_b[829] = 8'b11111111;
    mem_b[830] = 8'b00011111;
    mem_b[831] = 8'b00000000;
    mem_b[832] = 8'b00000000;
    mem_b[833] = 8'b11100000;
    mem_b[834] = 8'b11111111;
    mem_b[835] = 8'b11111111;
    mem_b[836] = 8'b11111111;
    mem_b[837] = 8'b11111111;
    mem_b[838] = 8'b11111111;
    mem_b[839] = 8'b11111111;
    mem_b[840] = 8'b11111111;
    mem_b[841] = 8'b11111111;
    mem_b[842] = 8'b11111111;
    mem_b[843] = 8'b11111111;
    mem_b[844] = 8'b11111111;
    mem_b[845] = 8'b11111111;
    mem_b[846] = 8'b00001111;
    mem_b[847] = 8'b00000000;
    mem_b[848] = 8'b00000000;
    mem_b[849] = 8'b11100000;
    mem_b[850] = 8'b11111111;
    mem_b[851] = 8'b11111111;
    mem_b[852] = 8'b11111111;
    mem_b[853] = 8'b11111111;
    mem_b[854] = 8'b11111111;
    mem_b[855] = 8'b11111111;
    mem_b[856] = 8'b11111111;
    mem_b[857] = 8'b11111111;
    mem_b[858] = 8'b11111111;
    mem_b[859] = 8'b11111111;
    mem_b[860] = 8'b11111111;
    mem_b[861] = 8'b11111111;
    mem_b[862] = 8'b00001111;
    mem_b[863] = 8'b00000000;
    mem_b[864] = 8'b00000000;
    mem_b[865] = 8'b11100000;
    mem_b[866] = 8'b11111111;
    mem_b[867] = 8'b11111111;
    mem_b[868] = 8'b11111111;
    mem_b[869] = 8'b11111111;
    mem_b[870] = 8'b11111111;
    mem_b[871] = 8'b11111111;
    mem_b[872] = 8'b11111111;
    mem_b[873] = 8'b11111111;
    mem_b[874] = 8'b11111111;
    mem_b[875] = 8'b11111111;
    mem_b[876] = 8'b11111111;
    mem_b[877] = 8'b11111111;
    mem_b[878] = 8'b00000111;
    mem_b[879] = 8'b00000000;
    mem_b[880] = 8'b00000000;
    mem_b[881] = 8'b11000000;
    mem_b[882] = 8'b11111111;
    mem_b[883] = 8'b11111111;
    mem_b[884] = 8'b11111111;
    mem_b[885] = 8'b11111111;
    mem_b[886] = 8'b11111111;
    mem_b[887] = 8'b11111111;
    mem_b[888] = 8'b11111111;
    mem_b[889] = 8'b11111111;
    mem_b[890] = 8'b11111111;
    mem_b[891] = 8'b11111111;
    mem_b[892] = 8'b11111111;
    mem_b[893] = 8'b11111111;
    mem_b[894] = 8'b00000011;
    mem_b[895] = 8'b00000000;
    mem_b[896] = 8'b00000000;
    mem_b[897] = 8'b11000000;
    mem_b[898] = 8'b11111111;
    mem_b[899] = 8'b11111111;
    mem_b[900] = 8'b11111111;
    mem_b[901] = 8'b11111111;
    mem_b[902] = 8'b11111111;
    mem_b[903] = 8'b11111111;
    mem_b[904] = 8'b11111111;
    mem_b[905] = 8'b11111111;
    mem_b[906] = 8'b11111111;
    mem_b[907] = 8'b11111111;
    mem_b[908] = 8'b11111111;
    mem_b[909] = 8'b11111111;
    mem_b[910] = 8'b00000001;
    mem_b[911] = 8'b00000000;
    mem_b[912] = 8'b00000000;
    mem_b[913] = 8'b10000000;
    mem_b[914] = 8'b11111111;
    mem_b[915] = 8'b11111111;
    mem_b[916] = 8'b11111111;
    mem_b[917] = 8'b11111111;
    mem_b[918] = 8'b11111111;
    mem_b[919] = 8'b11111111;
    mem_b[920] = 8'b11111111;
    mem_b[921] = 8'b11111111;
    mem_b[922] = 8'b11111111;
    mem_b[923] = 8'b11111111;
    mem_b[924] = 8'b11111111;
    mem_b[925] = 8'b11111111;
    mem_b[926] = 8'b00000000;
    mem_b[927] = 8'b00000000;
    mem_b[928] = 8'b00000000;
    mem_b[929] = 8'b10000000;
    mem_b[930] = 8'b11111111;
    mem_b[931] = 8'b11111111;
    mem_b[932] = 8'b11111111;
    mem_b[933] = 8'b11111111;
    mem_b[934] = 8'b11111111;
    mem_b[935] = 8'b11111111;
    mem_b[936] = 8'b11111111;
    mem_b[937] = 8'b11111111;
    mem_b[938] = 8'b11111111;
    mem_b[939] = 8'b11111111;
    mem_b[940] = 8'b11111111;
    mem_b[941] = 8'b11111111;
    mem_b[942] = 8'b11111111;
    mem_b[943] = 8'b00000111;
    mem_b[944] = 8'b00000000;
    mem_b[945] = 8'b10000000;
    mem_b[946] = 8'b11111111;
    mem_b[947] = 8'b11111111;
    mem_b[948] = 8'b11111111;
    mem_b[949] = 8'b11111111;
    mem_b[950] = 8'b11111111;
    mem_b[951] = 8'b11111111;
    mem_b[952] = 8'b11111111;
    mem_b[953] = 8'b11111111;
    mem_b[954] = 8'b11111111;
    mem_b[955] = 8'b11111111;
    mem_b[956] = 8'b11111111;
    mem_b[957] = 8'b11111111;
    mem_b[958] = 8'b11111111;
    mem_b[959] = 8'b00000111;
    mem_b[960] = 8'b00000000;
    mem_b[961] = 8'b00000000;
    mem_b[962] = 8'b11111111;
    mem_b[963] = 8'b11111111;
    mem_b[964] = 8'b11111111;
    mem_b[965] = 8'b11111111;
    mem_b[966] = 8'b11111111;
    mem_b[967] = 8'b11111111;
    mem_b[968] = 8'b11111111;
    mem_b[969] = 8'b11111111;
    mem_b[970] = 8'b11111111;
    mem_b[971] = 8'b11111111;
    mem_b[972] = 8'b11111111;
    mem_b[973] = 8'b11111111;
    mem_b[974] = 8'b11111111;
    mem_b[975] = 8'b00000111;
    mem_b[976] = 8'b11000000;
    mem_b[977] = 8'b00000001;
    mem_b[978] = 8'b11111111;
    mem_b[979] = 8'b11111111;
    mem_b[980] = 8'b11111111;
    mem_b[981] = 8'b11111111;
    mem_b[982] = 8'b11111111;
    mem_b[983] = 8'b11111111;
    mem_b[984] = 8'b11111111;
    mem_b[985] = 8'b11111111;
    mem_b[986] = 8'b11111111;
    mem_b[987] = 8'b11111111;
    mem_b[988] = 8'b11111111;
    mem_b[989] = 8'b11111111;
    mem_b[990] = 8'b11111111;
    mem_b[991] = 8'b00000111;
    mem_b[992] = 8'b11000000;
    mem_b[993] = 8'b00001111;
    mem_b[994] = 8'b11111110;
    mem_b[995] = 8'b11111111;
    mem_b[996] = 8'b11111111;
    mem_b[997] = 8'b11111111;
    mem_b[998] = 8'b11111111;
    mem_b[999] = 8'b11111111;
    mem_b[1000] = 8'b11111111;
    mem_b[1001] = 8'b11111111;
    mem_b[1002] = 8'b11111111;
    mem_b[1003] = 8'b11111111;
    mem_b[1004] = 8'b11111111;
    mem_b[1005] = 8'b11111111;
    mem_b[1006] = 8'b11111111;
    mem_b[1007] = 8'b00000011;
    mem_b[1008] = 8'b11000000;
    mem_b[1009] = 8'b11111111;
    mem_b[1010] = 8'b11111111;
    mem_b[1011] = 8'b11111111;
    mem_b[1012] = 8'b11111111;
    mem_b[1013] = 8'b11111111;
    mem_b[1014] = 8'b11111111;
    mem_b[1015] = 8'b11111111;
    mem_b[1016] = 8'b11111111;
    mem_b[1017] = 8'b11111111;
    mem_b[1018] = 8'b11111111;
    mem_b[1019] = 8'b11111111;
    mem_b[1020] = 8'b11111111;
    mem_b[1021] = 8'b11111111;
    mem_b[1022] = 8'b11111111;
    mem_b[1023] = 8'b00000001;
    mem_b[1024] = 8'b11000000;
    mem_b[1025] = 8'b11111111;
    mem_b[1026] = 8'b11111111;
    mem_b[1027] = 8'b11111111;
    mem_b[1028] = 8'b11111111;
    mem_b[1029] = 8'b11111111;
    mem_b[1030] = 8'b11111111;
    mem_b[1031] = 8'b11111111;
    mem_b[1032] = 8'b11111111;
    mem_b[1033] = 8'b11111111;
    mem_b[1034] = 8'b11111111;
    mem_b[1035] = 8'b11111111;
    mem_b[1036] = 8'b11111111;
    mem_b[1037] = 8'b11111111;
    mem_b[1038] = 8'b11111111;
    mem_b[1039] = 8'b00000001;
    mem_b[1040] = 8'b11000000;
    mem_b[1041] = 8'b11111111;
    mem_b[1042] = 8'b11111111;
    mem_b[1043] = 8'b11111111;
    mem_b[1044] = 8'b11111111;
    mem_b[1045] = 8'b11111111;
    mem_b[1046] = 8'b11111111;
    mem_b[1047] = 8'b11111111;
    mem_b[1048] = 8'b11111111;
    mem_b[1049] = 8'b11111111;
    mem_b[1050] = 8'b11111111;
    mem_b[1051] = 8'b11111111;
    mem_b[1052] = 8'b11111111;
    mem_b[1053] = 8'b11111111;
    mem_b[1054] = 8'b11111111;
    mem_b[1055] = 8'b00000000;
    mem_b[1056] = 8'b10000000;
    mem_b[1057] = 8'b11111111;
    mem_b[1058] = 8'b11111111;
    mem_b[1059] = 8'b11111111;
    mem_b[1060] = 8'b11111111;
    mem_b[1061] = 8'b11111111;
    mem_b[1062] = 8'b11111111;
    mem_b[1063] = 8'b11111111;
    mem_b[1064] = 8'b11111111;
    mem_b[1065] = 8'b11111111;
    mem_b[1066] = 8'b11111111;
    mem_b[1067] = 8'b11111111;
    mem_b[1068] = 8'b11111111;
    mem_b[1069] = 8'b11111111;
    mem_b[1070] = 8'b01111111;
    mem_b[1071] = 8'b00000000;
    mem_b[1072] = 8'b10000000;
    mem_b[1073] = 8'b11111111;
    mem_b[1074] = 8'b11111111;
    mem_b[1075] = 8'b11111111;
    mem_b[1076] = 8'b11111111;
    mem_b[1077] = 8'b11111111;
    mem_b[1078] = 8'b11111111;
    mem_b[1079] = 8'b11111111;
    mem_b[1080] = 8'b11111111;
    mem_b[1081] = 8'b11111111;
    mem_b[1082] = 8'b11111111;
    mem_b[1083] = 8'b11111111;
    mem_b[1084] = 8'b11111111;
    mem_b[1085] = 8'b11111111;
    mem_b[1086] = 8'b00111111;
    mem_b[1087] = 8'b00000000;
    mem_b[1088] = 8'b00000000;
    mem_b[1089] = 8'b11111111;
    mem_b[1090] = 8'b11111111;
    mem_b[1091] = 8'b11111111;
    mem_b[1092] = 8'b11111111;
    mem_b[1093] = 8'b11111111;
    mem_b[1094] = 8'b11111111;
    mem_b[1095] = 8'b11111111;
    mem_b[1096] = 8'b11111111;
    mem_b[1097] = 8'b11111111;
    mem_b[1098] = 8'b11111111;
    mem_b[1099] = 8'b11111111;
    mem_b[1100] = 8'b11111111;
    mem_b[1101] = 8'b01111111;
    mem_b[1102] = 8'b00011111;
    mem_b[1103] = 8'b00000000;
    mem_b[1104] = 8'b00000000;
    mem_b[1105] = 8'b11111110;
    mem_b[1106] = 8'b11111111;
    mem_b[1107] = 8'b11111111;
    mem_b[1108] = 8'b11111111;
    mem_b[1109] = 8'b11111111;
    mem_b[1110] = 8'b11111111;
    mem_b[1111] = 8'b11111111;
    mem_b[1112] = 8'b11111111;
    mem_b[1113] = 8'b11111111;
    mem_b[1114] = 8'b11111111;
    mem_b[1115] = 8'b11111111;
    mem_b[1116] = 8'b11111111;
    mem_b[1117] = 8'b11111111;
    mem_b[1118] = 8'b00011111;
    mem_b[1119] = 8'b00000000;
    mem_b[1120] = 8'b00000000;
    mem_b[1121] = 8'b11111110;
    mem_b[1122] = 8'b11111111;
    mem_b[1123] = 8'b11111111;
    mem_b[1124] = 8'b11111111;
    mem_b[1125] = 8'b11111111;
    mem_b[1126] = 8'b11111111;
    mem_b[1127] = 8'b11111111;
    mem_b[1128] = 8'b11111111;
    mem_b[1129] = 8'b11111111;
    mem_b[1130] = 8'b11111111;
    mem_b[1131] = 8'b11111111;
    mem_b[1132] = 8'b11111111;
    mem_b[1133] = 8'b11111111;
    mem_b[1134] = 8'b00001111;
    mem_b[1135] = 8'b00000000;
    mem_b[1136] = 8'b00000000;
    mem_b[1137] = 8'b11111100;
    mem_b[1138] = 8'b11111111;
    mem_b[1139] = 8'b11111111;
    mem_b[1140] = 8'b11111111;
    mem_b[1141] = 8'b11111111;
    mem_b[1142] = 8'b11111111;
    mem_b[1143] = 8'b11111111;
    mem_b[1144] = 8'b11111111;
    mem_b[1145] = 8'b11111111;
    mem_b[1146] = 8'b11111111;
    mem_b[1147] = 8'b11111111;
    mem_b[1148] = 8'b11111111;
    mem_b[1149] = 8'b11111111;
    mem_b[1150] = 8'b00000111;
    mem_b[1151] = 8'b00000000;
    mem_b[1152] = 8'b00000000;
    mem_b[1153] = 8'b11111000;
    mem_b[1154] = 8'b11111111;
    mem_b[1155] = 8'b11111111;
    mem_b[1156] = 8'b11111111;
    mem_b[1157] = 8'b11111111;
    mem_b[1158] = 8'b11111111;
    mem_b[1159] = 8'b11111111;
    mem_b[1160] = 8'b11111111;
    mem_b[1161] = 8'b11111111;
    mem_b[1162] = 8'b11111111;
    mem_b[1163] = 8'b11111111;
    mem_b[1164] = 8'b11111111;
    mem_b[1165] = 8'b11111111;
    mem_b[1166] = 8'b00000011;
    mem_b[1167] = 8'b00000000;
    mem_b[1168] = 8'b00000000;
    mem_b[1169] = 8'b11110000;
    mem_b[1170] = 8'b11111111;
    mem_b[1171] = 8'b11111111;
    mem_b[1172] = 8'b11111111;
    mem_b[1173] = 8'b11111111;
    mem_b[1174] = 8'b11111111;
    mem_b[1175] = 8'b11111111;
    mem_b[1176] = 8'b11111111;
    mem_b[1177] = 8'b11111111;
    mem_b[1178] = 8'b11111111;
    mem_b[1179] = 8'b11111111;
    mem_b[1180] = 8'b11111111;
    mem_b[1181] = 8'b11111111;
    mem_b[1182] = 8'b00000001;
    mem_b[1183] = 8'b00000000;
    mem_b[1184] = 8'b00000000;
    mem_b[1185] = 8'b11100000;
    mem_b[1186] = 8'b11111111;
    mem_b[1187] = 8'b11111111;
    mem_b[1188] = 8'b11111111;
    mem_b[1189] = 8'b11111111;
    mem_b[1190] = 8'b11111111;
    mem_b[1191] = 8'b11111111;
    mem_b[1192] = 8'b11111111;
    mem_b[1193] = 8'b11111111;
    mem_b[1194] = 8'b11111111;
    mem_b[1195] = 8'b11111111;
    mem_b[1196] = 8'b11111111;
    mem_b[1197] = 8'b11111111;
    mem_b[1198] = 8'b00000001;
    mem_b[1199] = 8'b00000000;
    mem_b[1200] = 8'b00000000;
    mem_b[1201] = 8'b11000000;
    mem_b[1202] = 8'b11111111;
    mem_b[1203] = 8'b11111111;
    mem_b[1204] = 8'b11111111;
    mem_b[1205] = 8'b11111111;
    mem_b[1206] = 8'b11111111;
    mem_b[1207] = 8'b11111111;
    mem_b[1208] = 8'b11111111;
    mem_b[1209] = 8'b11111111;
    mem_b[1210] = 8'b11111111;
    mem_b[1211] = 8'b11111111;
    mem_b[1212] = 8'b11111111;
    mem_b[1213] = 8'b11111111;
    mem_b[1214] = 8'b00000011;
    mem_b[1215] = 8'b00000000;
    mem_b[1216] = 8'b00000000;
    mem_b[1217] = 8'b10000000;
    mem_b[1218] = 8'b11111111;
    mem_b[1219] = 8'b11111111;
    mem_b[1220] = 8'b11111111;
    mem_b[1221] = 8'b11111111;
    mem_b[1222] = 8'b11111111;
    mem_b[1223] = 8'b11111111;
    mem_b[1224] = 8'b11111111;
    mem_b[1225] = 8'b11111111;
    mem_b[1226] = 8'b11111111;
    mem_b[1227] = 8'b11111111;
    mem_b[1228] = 8'b11111111;
    mem_b[1229] = 8'b11111111;
    mem_b[1230] = 8'b00000111;
    mem_b[1231] = 8'b00000000;
    mem_b[1232] = 8'b00000000;
    mem_b[1233] = 8'b11000000;
    mem_b[1234] = 8'b11111111;
    mem_b[1235] = 8'b11111111;
    mem_b[1236] = 8'b11111111;
    mem_b[1237] = 8'b11111111;
    mem_b[1238] = 8'b11111111;
    mem_b[1239] = 8'b11111111;
    mem_b[1240] = 8'b11111111;
    mem_b[1241] = 8'b11111111;
    mem_b[1242] = 8'b11111111;
    mem_b[1243] = 8'b11111111;
    mem_b[1244] = 8'b11111111;
    mem_b[1245] = 8'b11111111;
    mem_b[1246] = 8'b00001111;
    mem_b[1247] = 8'b00000000;
    mem_b[1248] = 8'b00000000;
    mem_b[1249] = 8'b11000000;
    mem_b[1250] = 8'b11111111;
    mem_b[1251] = 8'b11111111;
    mem_b[1252] = 8'b11111111;
    mem_b[1253] = 8'b11111111;
    mem_b[1254] = 8'b11111111;
    mem_b[1255] = 8'b11111111;
    mem_b[1256] = 8'b11111111;
    mem_b[1257] = 8'b11111111;
    mem_b[1258] = 8'b11111111;
    mem_b[1259] = 8'b11111111;
    mem_b[1260] = 8'b11111111;
    mem_b[1261] = 8'b11111111;
    mem_b[1262] = 8'b00001111;
    mem_b[1263] = 8'b00000000;
    mem_b[1264] = 8'b00000000;
    mem_b[1265] = 8'b11100000;
    mem_b[1266] = 8'b11111111;
    mem_b[1267] = 8'b11111111;
    mem_b[1268] = 8'b11111111;
    mem_b[1269] = 8'b11111111;
    mem_b[1270] = 8'b11111111;
    mem_b[1271] = 8'b11111111;
    mem_b[1272] = 8'b11111111;
    mem_b[1273] = 8'b11111111;
    mem_b[1274] = 8'b11111111;
    mem_b[1275] = 8'b11111111;
    mem_b[1276] = 8'b11111111;
    mem_b[1277] = 8'b11111111;
    mem_b[1278] = 8'b00011111;
    mem_b[1279] = 8'b00000000;
    mem_b[1280] = 8'b00000000;
    mem_b[1281] = 8'b11100000;
    mem_b[1282] = 8'b11111111;
    mem_b[1283] = 8'b11111111;
    mem_b[1284] = 8'b11111111;
    mem_b[1285] = 8'b11111111;
    mem_b[1286] = 8'b11111111;
    mem_b[1287] = 8'b11111111;
    mem_b[1288] = 8'b11111111;
    mem_b[1289] = 8'b11111111;
    mem_b[1290] = 8'b11111111;
    mem_b[1291] = 8'b11111111;
    mem_b[1292] = 8'b11111111;
    mem_b[1293] = 8'b11111111;
    mem_b[1294] = 8'b00111111;
    mem_b[1295] = 8'b00000000;
    mem_b[1296] = 8'b00000000;
    mem_b[1297] = 8'b11110000;
    mem_b[1298] = 8'b11111111;
    mem_b[1299] = 8'b11111111;
    mem_b[1300] = 8'b11111111;
    mem_b[1301] = 8'b11111111;
    mem_b[1302] = 8'b11111111;
    mem_b[1303] = 8'b11111111;
    mem_b[1304] = 8'b11111111;
    mem_b[1305] = 8'b11111111;
    mem_b[1306] = 8'b11111111;
    mem_b[1307] = 8'b11111111;
    mem_b[1308] = 8'b11111111;
    mem_b[1309] = 8'b11111111;
    mem_b[1310] = 8'b00111111;
    mem_b[1311] = 8'b00000000;
    mem_b[1312] = 8'b00000000;
    mem_b[1313] = 8'b11110000;
    mem_b[1314] = 8'b11111111;
    mem_b[1315] = 8'b11111111;
    mem_b[1316] = 8'b11111111;
    mem_b[1317] = 8'b11111111;
    mem_b[1318] = 8'b11111111;
    mem_b[1319] = 8'b11111111;
    mem_b[1320] = 8'b11111111;
    mem_b[1321] = 8'b11111111;
    mem_b[1322] = 8'b11111111;
    mem_b[1323] = 8'b11111111;
    mem_b[1324] = 8'b11111111;
    mem_b[1325] = 8'b11111111;
    mem_b[1326] = 8'b01111111;
    mem_b[1327] = 8'b00000000;
    mem_b[1328] = 8'b00000000;
    mem_b[1329] = 8'b11110000;
    mem_b[1330] = 8'b11111111;
    mem_b[1331] = 8'b11111111;
    mem_b[1332] = 8'b11111111;
    mem_b[1333] = 8'b11111111;
    mem_b[1334] = 8'b11111111;
    mem_b[1335] = 8'b11111111;
    mem_b[1336] = 8'b11111111;
    mem_b[1337] = 8'b11111111;
    mem_b[1338] = 8'b11111111;
    mem_b[1339] = 8'b11111111;
    mem_b[1340] = 8'b11111111;
    mem_b[1341] = 8'b11111111;
    mem_b[1342] = 8'b01111111;
    mem_b[1343] = 8'b00000000;
    mem_b[1344] = 8'b00000000;
    mem_b[1345] = 8'b11110000;
    mem_b[1346] = 8'b11111111;
    mem_b[1347] = 8'b11111111;
    mem_b[1348] = 8'b11111111;
    mem_b[1349] = 8'b11111111;
    mem_b[1350] = 8'b11111111;
    mem_b[1351] = 8'b11111111;
    mem_b[1352] = 8'b11111111;
    mem_b[1353] = 8'b11111111;
    mem_b[1354] = 8'b11111111;
    mem_b[1355] = 8'b11111111;
    mem_b[1356] = 8'b11111111;
    mem_b[1357] = 8'b11111111;
    mem_b[1358] = 8'b01111111;
    mem_b[1359] = 8'b00000000;
    mem_b[1360] = 8'b00000000;
    mem_b[1361] = 8'b11110000;
    mem_b[1362] = 8'b11111111;
    mem_b[1363] = 8'b11111111;
    mem_b[1364] = 8'b11111111;
    mem_b[1365] = 8'b11111111;
    mem_b[1366] = 8'b11111111;
    mem_b[1367] = 8'b11111111;
    mem_b[1368] = 8'b11111111;
    mem_b[1369] = 8'b11111111;
    mem_b[1370] = 8'b11111111;
    mem_b[1371] = 8'b11111111;
    mem_b[1372] = 8'b11111111;
    mem_b[1373] = 8'b11111111;
    mem_b[1374] = 8'b00111111;
    mem_b[1375] = 8'b00000000;
    mem_b[1376] = 8'b00000000;
    mem_b[1377] = 8'b11110000;
    mem_b[1378] = 8'b11111111;
    mem_b[1379] = 8'b11111111;
    mem_b[1380] = 8'b11111111;
    mem_b[1381] = 8'b11111111;
    mem_b[1382] = 8'b11111111;
    mem_b[1383] = 8'b11111111;
    mem_b[1384] = 8'b11111111;
    mem_b[1385] = 8'b11111111;
    mem_b[1386] = 8'b11111111;
    mem_b[1387] = 8'b11111111;
    mem_b[1388] = 8'b11111111;
    mem_b[1389] = 8'b11111111;
    mem_b[1390] = 8'b00011111;
    mem_b[1391] = 8'b00000000;
    mem_b[1392] = 8'b00000000;
    mem_b[1393] = 8'b11110000;
    mem_b[1394] = 8'b11111111;
    mem_b[1395] = 8'b11111111;
    mem_b[1396] = 8'b11111111;
    mem_b[1397] = 8'b11111111;
    mem_b[1398] = 8'b11111111;
    mem_b[1399] = 8'b11111111;
    mem_b[1400] = 8'b11111111;
    mem_b[1401] = 8'b11111111;
    mem_b[1402] = 8'b11111111;
    mem_b[1403] = 8'b11111111;
    mem_b[1404] = 8'b11111111;
    mem_b[1405] = 8'b11111111;
    mem_b[1406] = 8'b00000111;
    mem_b[1407] = 8'b00000000;
    mem_b[1408] = 8'b00000000;
    mem_b[1409] = 8'b11110000;
    mem_b[1410] = 8'b11111111;
    mem_b[1411] = 8'b11111111;
    mem_b[1412] = 8'b11111111;
    mem_b[1413] = 8'b11111111;
    mem_b[1414] = 8'b11111111;
    mem_b[1415] = 8'b11111111;
    mem_b[1416] = 8'b11111111;
    mem_b[1417] = 8'b11111111;
    mem_b[1418] = 8'b11111111;
    mem_b[1419] = 8'b11111111;
    mem_b[1420] = 8'b11110111;
    mem_b[1421] = 8'b11111111;
    mem_b[1422] = 8'b00000000;
    mem_b[1423] = 8'b00000000;
    mem_b[1424] = 8'b00000000;
    mem_b[1425] = 8'b11110000;
    mem_b[1426] = 8'b11111111;
    mem_b[1427] = 8'b11111111;
    mem_b[1428] = 8'b11111111;
    mem_b[1429] = 8'b11111111;
    mem_b[1430] = 8'b11111111;
    mem_b[1431] = 8'b11111111;
    mem_b[1432] = 8'b11111111;
    mem_b[1433] = 8'b11111111;
    mem_b[1434] = 8'b11111111;
    mem_b[1435] = 8'b11111111;
    mem_b[1436] = 8'b11110011;
    mem_b[1437] = 8'b00000111;
    mem_b[1438] = 8'b00000000;
    mem_b[1439] = 8'b00000000;
    mem_b[1440] = 8'b00000000;
    mem_b[1441] = 8'b10000000;
    mem_b[1442] = 8'b11111111;
    mem_b[1443] = 8'b11110011;
    mem_b[1444] = 8'b11111111;
    mem_b[1445] = 8'b11111111;
    mem_b[1446] = 8'b11111111;
    mem_b[1447] = 8'b11111111;
    mem_b[1448] = 8'b11111111;
    mem_b[1449] = 8'b11111111;
    mem_b[1450] = 8'b11111111;
    mem_b[1451] = 8'b11111111;
    mem_b[1452] = 8'b00000001;
    mem_b[1453] = 8'b00000000;
    mem_b[1454] = 8'b00000000;
    mem_b[1455] = 8'b00000000;
    mem_b[1456] = 8'b00000000;
    mem_b[1457] = 8'b00000000;
    mem_b[1458] = 8'b00000000;
    mem_b[1459] = 8'b11000000;
    mem_b[1460] = 8'b11111111;
    mem_b[1461] = 8'b11111111;
    mem_b[1462] = 8'b11111111;
    mem_b[1463] = 8'b11111111;
    mem_b[1464] = 8'b11111111;
    mem_b[1465] = 8'b11111111;
    mem_b[1466] = 8'b11111111;
    mem_b[1467] = 8'b01111111;
    mem_b[1468] = 8'b00000000;
    mem_b[1469] = 8'b00000000;
    mem_b[1470] = 8'b00000000;
    mem_b[1471] = 8'b00000000;
    mem_b[1472] = 8'b00000000;
    mem_b[1473] = 8'b00000000;
    mem_b[1474] = 8'b00000000;
    mem_b[1475] = 8'b10000000;
    mem_b[1476] = 8'b11111111;
    mem_b[1477] = 8'b11111111;
    mem_b[1478] = 8'b11111111;
    mem_b[1479] = 8'b11111111;
    mem_b[1480] = 8'b11111111;
    mem_b[1481] = 8'b11111111;
    mem_b[1482] = 8'b11111111;
    mem_b[1483] = 8'b00011111;
    mem_b[1484] = 8'b00000000;
    mem_b[1485] = 8'b00000000;
    mem_b[1486] = 8'b00000000;
    mem_b[1487] = 8'b00000000;
    mem_b[1488] = 8'b00000000;
    mem_b[1489] = 8'b00000000;
    mem_b[1490] = 8'b00000000;
    mem_b[1491] = 8'b00000000;
    mem_b[1492] = 8'b11111110;
    mem_b[1493] = 8'b11111111;
    mem_b[1494] = 8'b11111111;
    mem_b[1495] = 8'b11111111;
    mem_b[1496] = 8'b11111111;
    mem_b[1497] = 8'b11111111;
    mem_b[1498] = 8'b11111111;
    mem_b[1499] = 8'b00000011;
    mem_b[1500] = 8'b00000000;
    mem_b[1501] = 8'b00000000;
    mem_b[1502] = 8'b00000000;
    mem_b[1503] = 8'b00000000;
    mem_b[1504] = 8'b00000000;
    mem_b[1505] = 8'b00000000;
    mem_b[1506] = 8'b00000000;
    mem_b[1507] = 8'b00000000;
    mem_b[1508] = 8'b11111000;
    mem_b[1509] = 8'b11111111;
    mem_b[1510] = 8'b11111111;
    mem_b[1511] = 8'b11111111;
    mem_b[1512] = 8'b11111111;
    mem_b[1513] = 8'b11111111;
    mem_b[1514] = 8'b11111111;
    mem_b[1515] = 8'b00000001;
    mem_b[1516] = 8'b00000000;
    mem_b[1517] = 8'b00000000;
    mem_b[1518] = 8'b00000000;
    mem_b[1519] = 8'b00000000;
    mem_b[1520] = 8'b00000000;
    mem_b[1521] = 8'b00000000;
    mem_b[1522] = 8'b00000000;
    mem_b[1523] = 8'b00000000;
    mem_b[1524] = 8'b11100000;
    mem_b[1525] = 8'b11111111;
    mem_b[1526] = 8'b11111111;
    mem_b[1527] = 8'b11111111;
    mem_b[1528] = 8'b11111111;
    mem_b[1529] = 8'b11111111;
    mem_b[1530] = 8'b11111111;
    mem_b[1531] = 8'b00000001;
    mem_b[1532] = 8'b00000000;
    mem_b[1533] = 8'b00000000;
    mem_b[1534] = 8'b00000000;
    mem_b[1535] = 8'b00000000;
    mem_b[1536] = 8'b00000000;
    mem_b[1537] = 8'b00000000;
    mem_b[1538] = 8'b00000000;
    mem_b[1539] = 8'b00000000;
    mem_b[1540] = 8'b11100000;
    mem_b[1541] = 8'b11111111;
    mem_b[1542] = 8'b11111111;
    mem_b[1543] = 8'b11111111;
    mem_b[1544] = 8'b11111111;
    mem_b[1545] = 8'b11111111;
    mem_b[1546] = 8'b11111111;
    mem_b[1547] = 8'b00000011;
    mem_b[1548] = 8'b00000000;
    mem_b[1549] = 8'b00000000;
    mem_b[1550] = 8'b00000000;
    mem_b[1551] = 8'b00000000;
    mem_b[1552] = 8'b00000000;
    mem_b[1553] = 8'b00000000;
    mem_b[1554] = 8'b00000000;
    mem_b[1555] = 8'b00000000;
    mem_b[1556] = 8'b11000000;
    mem_b[1557] = 8'b11111111;
    mem_b[1558] = 8'b11111111;
    mem_b[1559] = 8'b11111111;
    mem_b[1560] = 8'b11111111;
    mem_b[1561] = 8'b11111111;
    mem_b[1562] = 8'b11111111;
    mem_b[1563] = 8'b00000011;
    mem_b[1564] = 8'b00000000;
    mem_b[1565] = 8'b00000000;
    mem_b[1566] = 8'b00000000;
    mem_b[1567] = 8'b00000000;
    mem_b[1568] = 8'b00000000;
    mem_b[1569] = 8'b00000000;
    mem_b[1570] = 8'b00000000;
    mem_b[1571] = 8'b00000000;
    mem_b[1572] = 8'b11000000;
    mem_b[1573] = 8'b11111111;
    mem_b[1574] = 8'b11111111;
    mem_b[1575] = 8'b11111111;
    mem_b[1576] = 8'b11111111;
    mem_b[1577] = 8'b11111111;
    mem_b[1578] = 8'b11111111;
    mem_b[1579] = 8'b00000111;
    mem_b[1580] = 8'b00000000;
    mem_b[1581] = 8'b00000000;
    mem_b[1582] = 8'b00000000;
    mem_b[1583] = 8'b00000000;
    mem_b[1584] = 8'b00000000;
    mem_b[1585] = 8'b00000000;
    mem_b[1586] = 8'b00000000;
    mem_b[1587] = 8'b00000000;
    mem_b[1588] = 8'b10000000;
    mem_b[1589] = 8'b11111111;
    mem_b[1590] = 8'b11111111;
    mem_b[1591] = 8'b11111111;
    mem_b[1592] = 8'b11111111;
    mem_b[1593] = 8'b11111111;
    mem_b[1594] = 8'b11111111;
    mem_b[1595] = 8'b00001111;
    mem_b[1596] = 8'b00000000;
    mem_b[1597] = 8'b00000000;
    mem_b[1598] = 8'b00000000;
    mem_b[1599] = 8'b00000000;
    mem_b[1600] = 8'b00000000;
    mem_b[1601] = 8'b00000000;
    mem_b[1602] = 8'b00000000;
    mem_b[1603] = 8'b00000000;
    mem_b[1604] = 8'b10000000;
    mem_b[1605] = 8'b11111111;
    mem_b[1606] = 8'b11111111;
    mem_b[1607] = 8'b11111111;
    mem_b[1608] = 8'b11111111;
    mem_b[1609] = 8'b11111111;
    mem_b[1610] = 8'b11111111;
    mem_b[1611] = 8'b00001111;
    mem_b[1612] = 8'b00000000;
    mem_b[1613] = 8'b00000000;
    mem_b[1614] = 8'b00000000;
    mem_b[1615] = 8'b00000000;
    mem_b[1616] = 8'b00000000;
    mem_b[1617] = 8'b00000000;
    mem_b[1618] = 8'b00000000;
    mem_b[1619] = 8'b00000000;
    mem_b[1620] = 8'b00000000;
    mem_b[1621] = 8'b11111111;
    mem_b[1622] = 8'b11111111;
    mem_b[1623] = 8'b11111111;
    mem_b[1624] = 8'b11111111;
    mem_b[1625] = 8'b11111111;
    mem_b[1626] = 8'b11111111;
    mem_b[1627] = 8'b00001111;
    mem_b[1628] = 8'b00000000;
    mem_b[1629] = 8'b00000000;
    mem_b[1630] = 8'b00000000;
    mem_b[1631] = 8'b00000000;
    mem_b[1632] = 8'b00000000;
    mem_b[1633] = 8'b00000000;
    mem_b[1634] = 8'b00000000;
    mem_b[1635] = 8'b00000000;
    mem_b[1636] = 8'b00000000;
    mem_b[1637] = 8'b11111110;
    mem_b[1638] = 8'b11111111;
    mem_b[1639] = 8'b11111111;
    mem_b[1640] = 8'b11111111;
    mem_b[1641] = 8'b11111111;
    mem_b[1642] = 8'b11111111;
    mem_b[1643] = 8'b00011111;
    mem_b[1644] = 8'b00000000;
    mem_b[1645] = 8'b00000000;
    mem_b[1646] = 8'b00000000;
    mem_b[1647] = 8'b00000000;
    mem_b[1648] = 8'b00000000;
    mem_b[1649] = 8'b00000000;
    mem_b[1650] = 8'b00000000;
    mem_b[1651] = 8'b00000000;
    mem_b[1652] = 8'b00000000;
    mem_b[1653] = 8'b11111100;
    mem_b[1654] = 8'b11111111;
    mem_b[1655] = 8'b11111111;
    mem_b[1656] = 8'b11111111;
    mem_b[1657] = 8'b11111111;
    mem_b[1658] = 8'b11111111;
    mem_b[1659] = 8'b00011111;
    mem_b[1660] = 8'b00000000;
    mem_b[1661] = 8'b00000000;
    mem_b[1662] = 8'b00000000;
    mem_b[1663] = 8'b00000000;
    mem_b[1664] = 8'b00000000;
    mem_b[1665] = 8'b00000000;
    mem_b[1666] = 8'b00000000;
    mem_b[1667] = 8'b00000000;
    mem_b[1668] = 8'b00000000;
    mem_b[1669] = 8'b11111000;
    mem_b[1670] = 8'b11111111;
    mem_b[1671] = 8'b11111111;
    mem_b[1672] = 8'b11111111;
    mem_b[1673] = 8'b11111111;
    mem_b[1674] = 8'b11111111;
    mem_b[1675] = 8'b00111111;
    mem_b[1676] = 8'b00000000;
    mem_b[1677] = 8'b00000000;
    mem_b[1678] = 8'b00000000;
    mem_b[1679] = 8'b00000000;
    mem_b[1680] = 8'b00000000;
    mem_b[1681] = 8'b00000000;
    mem_b[1682] = 8'b00000000;
    mem_b[1683] = 8'b00000000;
    mem_b[1684] = 8'b00000000;
    mem_b[1685] = 8'b11111100;
    mem_b[1686] = 8'b11111111;
    mem_b[1687] = 8'b11111111;
    mem_b[1688] = 8'b11111111;
    mem_b[1689] = 8'b11111111;
    mem_b[1690] = 8'b11111111;
    mem_b[1691] = 8'b00111111;
    mem_b[1692] = 8'b00000000;
    mem_b[1693] = 8'b00000000;
    mem_b[1694] = 8'b00000000;
    mem_b[1695] = 8'b00000000;
    mem_b[1696] = 8'b00000000;
    mem_b[1697] = 8'b00000000;
    mem_b[1698] = 8'b00000000;
    mem_b[1699] = 8'b00000000;
    mem_b[1700] = 8'b00000000;
    mem_b[1701] = 8'b11111100;
    mem_b[1702] = 8'b11111111;
    mem_b[1703] = 8'b11111111;
    mem_b[1704] = 8'b11111111;
    mem_b[1705] = 8'b11111111;
    mem_b[1706] = 8'b11111111;
    mem_b[1707] = 8'b00111111;
    mem_b[1708] = 8'b00000000;
    mem_b[1709] = 8'b00000000;
    mem_b[1710] = 8'b00000000;
    mem_b[1711] = 8'b00000000;
    mem_b[1712] = 8'b00000000;
    mem_b[1713] = 8'b00000000;
    mem_b[1714] = 8'b00000000;
    mem_b[1715] = 8'b00000000;
    mem_b[1716] = 8'b00000000;
    mem_b[1717] = 8'b11111110;
    mem_b[1718] = 8'b11111111;
    mem_b[1719] = 8'b11111111;
    mem_b[1720] = 8'b11111111;
    mem_b[1721] = 8'b11111111;
    mem_b[1722] = 8'b11111111;
    mem_b[1723] = 8'b00111111;
    mem_b[1724] = 8'b00000000;
    mem_b[1725] = 8'b00000000;
    mem_b[1726] = 8'b00000000;
    mem_b[1727] = 8'b00000000;
    mem_b[1728] = 8'b00000000;
    mem_b[1729] = 8'b00000000;
    mem_b[1730] = 8'b00000000;
    mem_b[1731] = 8'b00000000;
    mem_b[1732] = 8'b00000000;
    mem_b[1733] = 8'b11111111;
    mem_b[1734] = 8'b11111111;
    mem_b[1735] = 8'b11111111;
    mem_b[1736] = 8'b11111111;
    mem_b[1737] = 8'b11111111;
    mem_b[1738] = 8'b11111111;
    mem_b[1739] = 8'b01111111;
    mem_b[1740] = 8'b00000000;
    mem_b[1741] = 8'b00000000;
    mem_b[1742] = 8'b00000000;
    mem_b[1743] = 8'b00000000;
    mem_b[1744] = 8'b00000000;
    mem_b[1745] = 8'b00000000;
    mem_b[1746] = 8'b00000000;
    mem_b[1747] = 8'b00000000;
    mem_b[1748] = 8'b10000000;
    mem_b[1749] = 8'b11111111;
    mem_b[1750] = 8'b11111111;
    mem_b[1751] = 8'b11111111;
    mem_b[1752] = 8'b11111111;
    mem_b[1753] = 8'b11111111;
    mem_b[1754] = 8'b11111111;
    mem_b[1755] = 8'b01111111;
    mem_b[1756] = 8'b00000000;
    mem_b[1757] = 8'b00000000;
    mem_b[1758] = 8'b00000000;
    mem_b[1759] = 8'b00000000;
    mem_b[1760] = 8'b00000000;
    mem_b[1761] = 8'b00000000;
    mem_b[1762] = 8'b00000000;
    mem_b[1763] = 8'b00000000;
    mem_b[1764] = 8'b11000000;
    mem_b[1765] = 8'b11111111;
    mem_b[1766] = 8'b11111111;
    mem_b[1767] = 8'b11111111;
    mem_b[1768] = 8'b11111111;
    mem_b[1769] = 8'b11111111;
    mem_b[1770] = 8'b11111111;
    mem_b[1771] = 8'b01111111;
    mem_b[1772] = 8'b00000000;
    mem_b[1773] = 8'b00000000;
    mem_b[1774] = 8'b00000000;
    mem_b[1775] = 8'b00000000;
    mem_b[1776] = 8'b00000000;
    mem_b[1777] = 8'b00000000;
    mem_b[1778] = 8'b00000000;
    mem_b[1779] = 8'b00000000;
    mem_b[1780] = 8'b11000000;
    mem_b[1781] = 8'b11111111;
    mem_b[1782] = 8'b11111111;
    mem_b[1783] = 8'b11111111;
    mem_b[1784] = 8'b11111111;
    mem_b[1785] = 8'b11111111;
    mem_b[1786] = 8'b11111111;
    mem_b[1787] = 8'b11111111;
    mem_b[1788] = 8'b00000000;
    mem_b[1789] = 8'b00000000;
    mem_b[1790] = 8'b00000000;
    mem_b[1791] = 8'b00000000;
    mem_b[1792] = 8'b00000000;
    mem_b[1793] = 8'b00000000;
    mem_b[1794] = 8'b00000000;
    mem_b[1795] = 8'b00000000;
    mem_b[1796] = 8'b11000000;
    mem_b[1797] = 8'b11111111;
    mem_b[1798] = 8'b11111111;
    mem_b[1799] = 8'b11111111;
    mem_b[1800] = 8'b11111111;
    mem_b[1801] = 8'b11111111;
    mem_b[1802] = 8'b11111111;
    mem_b[1803] = 8'b11111111;
    mem_b[1804] = 8'b00000000;
    mem_b[1805] = 8'b00000000;
    mem_b[1806] = 8'b00000000;
    mem_b[1807] = 8'b00000000;
    mem_b[1808] = 8'b00000000;
    mem_b[1809] = 8'b00000000;
    mem_b[1810] = 8'b00000000;
    mem_b[1811] = 8'b00000000;
    mem_b[1812] = 8'b11000000;
    mem_b[1813] = 8'b11111111;
    mem_b[1814] = 8'b11111111;
    mem_b[1815] = 8'b11111111;
    mem_b[1816] = 8'b11111111;
    mem_b[1817] = 8'b11111111;
    mem_b[1818] = 8'b11111111;
    mem_b[1819] = 8'b11111111;
    mem_b[1820] = 8'b00000000;
    mem_b[1821] = 8'b00000000;
    mem_b[1822] = 8'b00000000;
    mem_b[1823] = 8'b00000000;
    mem_b[1824] = 8'b00000000;
    mem_b[1825] = 8'b00000000;
    mem_b[1826] = 8'b00000000;
    mem_b[1827] = 8'b00000000;
    mem_b[1828] = 8'b00000000;
    mem_b[1829] = 8'b11100000;
    mem_b[1830] = 8'b11111111;
    mem_b[1831] = 8'b11111111;
    mem_b[1832] = 8'b11111111;
    mem_b[1833] = 8'b11111111;
    mem_b[1834] = 8'b11111111;
    mem_b[1835] = 8'b11111111;
    mem_b[1836] = 8'b00000000;
    mem_b[1837] = 8'b00000000;
    mem_b[1838] = 8'b00000000;
    mem_b[1839] = 8'b00000000;
    mem_b[1840] = 8'b00000000;
    mem_b[1841] = 8'b00000000;
    mem_b[1842] = 8'b00000000;
    mem_b[1843] = 8'b00000000;
    mem_b[1844] = 8'b00000000;
    mem_b[1845] = 8'b11100000;
    mem_b[1846] = 8'b11111111;
    mem_b[1847] = 8'b11111111;
    mem_b[1848] = 8'b11111111;
    mem_b[1849] = 8'b11111111;
    mem_b[1850] = 8'b11111111;
    mem_b[1851] = 8'b11111111;
    mem_b[1852] = 8'b00000001;
    mem_b[1853] = 8'b00000000;
    mem_b[1854] = 8'b00000000;
    mem_b[1855] = 8'b00000000;
    mem_b[1856] = 8'b00000000;
    mem_b[1857] = 8'b00000000;
    mem_b[1858] = 8'b00000000;
    mem_b[1859] = 8'b00000000;
    mem_b[1860] = 8'b00000000;
    mem_b[1861] = 8'b11100000;
    mem_b[1862] = 8'b11111111;
    mem_b[1863] = 8'b11111111;
    mem_b[1864] = 8'b11111111;
    mem_b[1865] = 8'b11111111;
    mem_b[1866] = 8'b11111111;
    mem_b[1867] = 8'b11111111;
    mem_b[1868] = 8'b00000001;
    mem_b[1869] = 8'b00000000;
    mem_b[1870] = 8'b00000000;
    mem_b[1871] = 8'b00000000;
    mem_b[1872] = 8'b00000000;
    mem_b[1873] = 8'b00000000;
    mem_b[1874] = 8'b00000000;
    mem_b[1875] = 8'b00000000;
    mem_b[1876] = 8'b00000000;
    mem_b[1877] = 8'b11110000;
    mem_b[1878] = 8'b11111111;
    mem_b[1879] = 8'b11111111;
    mem_b[1880] = 8'b11111111;
    mem_b[1881] = 8'b11111111;
    mem_b[1882] = 8'b11111111;
    mem_b[1883] = 8'b11111111;
    mem_b[1884] = 8'b00000001;
    mem_b[1885] = 8'b00000000;
    mem_b[1886] = 8'b00000000;
    mem_b[1887] = 8'b00000000;
    mem_b[1888] = 8'b00000000;
    mem_b[1889] = 8'b00000000;
    mem_b[1890] = 8'b00000000;
    mem_b[1891] = 8'b00000000;
    mem_b[1892] = 8'b00000000;
    mem_b[1893] = 8'b11110000;
    mem_b[1894] = 8'b11111111;
    mem_b[1895] = 8'b11111111;
    mem_b[1896] = 8'b11111111;
    mem_b[1897] = 8'b11111111;
    mem_b[1898] = 8'b11111111;
    mem_b[1899] = 8'b11111111;
    mem_b[1900] = 8'b00000001;
    mem_b[1901] = 8'b00000000;
    mem_b[1902] = 8'b00000000;
    mem_b[1903] = 8'b00000000;
    mem_b[1904] = 8'b00000000;
    mem_b[1905] = 8'b00000000;
    mem_b[1906] = 8'b00000000;
    mem_b[1907] = 8'b00000000;
    mem_b[1908] = 8'b00000000;
    mem_b[1909] = 8'b11110000;
    mem_b[1910] = 8'b11111111;
    mem_b[1911] = 8'b11111111;
    mem_b[1912] = 8'b11111111;
    mem_b[1913] = 8'b11111111;
    mem_b[1914] = 8'b11111111;
    mem_b[1915] = 8'b11111111;
    mem_b[1916] = 8'b00000011;
    mem_b[1917] = 8'b00000000;
    mem_b[1918] = 8'b00000000;
    mem_b[1919] = 8'b00000000;
    mem_b[1920] = 8'b00000000;
    mem_b[1921] = 8'b00000000;
    mem_b[1922] = 8'b00000000;
    mem_b[1923] = 8'b00000000;
    mem_b[1924] = 8'b00000000;
    mem_b[1925] = 8'b11111000;
    mem_b[1926] = 8'b11111111;
    mem_b[1927] = 8'b11111111;
    mem_b[1928] = 8'b11111111;
    mem_b[1929] = 8'b11111111;
    mem_b[1930] = 8'b11111111;
    mem_b[1931] = 8'b11111111;
    mem_b[1932] = 8'b00000011;
    mem_b[1933] = 8'b00000000;
    mem_b[1934] = 8'b00000000;
    mem_b[1935] = 8'b00000000;
    mem_b[1936] = 8'b00000000;
    mem_b[1937] = 8'b00000000;
    mem_b[1938] = 8'b00000000;
    mem_b[1939] = 8'b00000000;
    mem_b[1940] = 8'b00000000;
    mem_b[1941] = 8'b11111000;
    mem_b[1942] = 8'b11111111;
    mem_b[1943] = 8'b11111111;
    mem_b[1944] = 8'b11111111;
    mem_b[1945] = 8'b11111111;
    mem_b[1946] = 8'b11111111;
    mem_b[1947] = 8'b11111111;
    mem_b[1948] = 8'b00000011;
    mem_b[1949] = 8'b00000000;
    mem_b[1950] = 8'b00000000;
    mem_b[1951] = 8'b00000000;
    mem_b[1952] = 8'b00000000;
    mem_b[1953] = 8'b00000000;
    mem_b[1954] = 8'b00000000;
    mem_b[1955] = 8'b00000000;
    mem_b[1956] = 8'b00000000;
    mem_b[1957] = 8'b11111000;
    mem_b[1958] = 8'b11111111;
    mem_b[1959] = 8'b11111111;
    mem_b[1960] = 8'b11111111;
    mem_b[1961] = 8'b11111111;
    mem_b[1962] = 8'b11111111;
    mem_b[1963] = 8'b11111111;
    mem_b[1964] = 8'b00000011;
    mem_b[1965] = 8'b00000000;
    mem_b[1966] = 8'b00000000;
    mem_b[1967] = 8'b00000000;
    mem_b[1968] = 8'b00000000;
    mem_b[1969] = 8'b00000000;
    mem_b[1970] = 8'b00000000;
    mem_b[1971] = 8'b00000000;
    mem_b[1972] = 8'b00000000;
    mem_b[1973] = 8'b11111000;
    mem_b[1974] = 8'b11111111;
    mem_b[1975] = 8'b11111111;
    mem_b[1976] = 8'b11111111;
    mem_b[1977] = 8'b11111111;
    mem_b[1978] = 8'b11111111;
    mem_b[1979] = 8'b11111111;
    mem_b[1980] = 8'b00000011;
    mem_b[1981] = 8'b00000000;
    mem_b[1982] = 8'b00000000;
    mem_b[1983] = 8'b00000000;
    mem_b[1984] = 8'b00000000;
    mem_b[1985] = 8'b00000000;
    mem_b[1986] = 8'b00000000;
    mem_b[1987] = 8'b00000000;
    mem_b[1988] = 8'b00000000;
    mem_b[1989] = 8'b11111000;
    mem_b[1990] = 8'b11111111;
    mem_b[1991] = 8'b11111111;
    mem_b[1992] = 8'b11111111;
    mem_b[1993] = 8'b11111111;
    mem_b[1994] = 8'b11111111;
    mem_b[1995] = 8'b11111111;
    mem_b[1996] = 8'b00000011;
    mem_b[1997] = 8'b00000000;
    mem_b[1998] = 8'b00000000;
    mem_b[1999] = 8'b00000000;
    mem_b[2000] = 8'b00000000;
    mem_b[2001] = 8'b00000000;
    mem_b[2002] = 8'b00000000;
    mem_b[2003] = 8'b00000000;
    mem_b[2004] = 8'b00000000;
    mem_b[2005] = 8'b11111000;
    mem_b[2006] = 8'b11111111;
    mem_b[2007] = 8'b11111111;
    mem_b[2008] = 8'b11111111;
    mem_b[2009] = 8'b11111111;
    mem_b[2010] = 8'b11111111;
    mem_b[2011] = 8'b11111111;
    mem_b[2012] = 8'b00000011;
    mem_b[2013] = 8'b00000000;
    mem_b[2014] = 8'b00000000;
    mem_b[2015] = 8'b00000000;
    mem_b[2016] = 8'b00000000;
    mem_b[2017] = 8'b00000000;
    mem_b[2018] = 8'b00000000;
    mem_b[2019] = 8'b00000000;
    mem_b[2020] = 8'b00000000;
    mem_b[2021] = 8'b11111000;
    mem_b[2022] = 8'b11111111;
    mem_b[2023] = 8'b11111111;
    mem_b[2024] = 8'b11111111;
    mem_b[2025] = 8'b11111111;
    mem_b[2026] = 8'b11111111;
    mem_b[2027] = 8'b11111111;
    mem_b[2028] = 8'b00000011;
    mem_b[2029] = 8'b00000000;
    mem_b[2030] = 8'b00000000;
    mem_b[2031] = 8'b00000000;
    mem_b[2032] = 8'b00000000;
    mem_b[2033] = 8'b00000000;
    mem_b[2034] = 8'b00000000;
    mem_b[2035] = 8'b00000000;
    mem_b[2036] = 8'b00000000;
    mem_b[2037] = 8'b11111000;
    mem_b[2038] = 8'b11111111;
    mem_b[2039] = 8'b11111111;
    mem_b[2040] = 8'b11111111;
    mem_b[2041] = 8'b11111111;
    mem_b[2042] = 8'b11111111;
    mem_b[2043] = 8'b11111111;
    mem_b[2044] = 8'b00000011;
    mem_b[2045] = 8'b00000000;
    mem_b[2046] = 8'b00000000;
    mem_b[2047] = 8'b00000000;
end

reg [7:0] mem_c [0:2047];
initial begin
    mem_c[0] = 8'b00000000;
    mem_c[1] = 8'b00000000;
    mem_c[2] = 8'b00000000;
    mem_c[3] = 8'b00000000;
    mem_c[4] = 8'b00000000;
    mem_c[5] = 8'b00000000;
    mem_c[6] = 8'b00000000;
    mem_c[7] = 8'b00000000;
    mem_c[8] = 8'b00000000;
    mem_c[9] = 8'b00000000;
    mem_c[10] = 8'b00000000;
    mem_c[11] = 8'b00000000;
    mem_c[12] = 8'b00000000;
    mem_c[13] = 8'b00000000;
    mem_c[14] = 8'b00000000;
    mem_c[15] = 8'b00000000;
    mem_c[16] = 8'b00000000;
    mem_c[17] = 8'b00000000;
    mem_c[18] = 8'b00000000;
    mem_c[19] = 8'b00000000;
    mem_c[20] = 8'b00000000;
    mem_c[21] = 8'b00000000;
    mem_c[22] = 8'b00000000;
    mem_c[23] = 8'b00000000;
    mem_c[24] = 8'b00000000;
    mem_c[25] = 8'b00000000;
    mem_c[26] = 8'b00000000;
    mem_c[27] = 8'b00000000;
    mem_c[28] = 8'b00000000;
    mem_c[29] = 8'b00000000;
    mem_c[30] = 8'b00000000;
    mem_c[31] = 8'b00000000;
    mem_c[32] = 8'b00000000;
    mem_c[33] = 8'b00000000;
    mem_c[34] = 8'b00000000;
    mem_c[35] = 8'b00000000;
    mem_c[36] = 8'b00000000;
    mem_c[37] = 8'b00000000;
    mem_c[38] = 8'b00000000;
    mem_c[39] = 8'b00000000;
    mem_c[40] = 8'b00000000;
    mem_c[41] = 8'b00000000;
    mem_c[42] = 8'b00000000;
    mem_c[43] = 8'b00000000;
    mem_c[44] = 8'b00000000;
    mem_c[45] = 8'b00000000;
    mem_c[46] = 8'b00000000;
    mem_c[47] = 8'b00000000;
    mem_c[48] = 8'b00000000;
    mem_c[49] = 8'b00000000;
    mem_c[50] = 8'b00000000;
    mem_c[51] = 8'b00000000;
    mem_c[52] = 8'b00000000;
    mem_c[53] = 8'b00000000;
    mem_c[54] = 8'b00000000;
    mem_c[55] = 8'b00000000;
    mem_c[56] = 8'b00000000;
    mem_c[57] = 8'b00000000;
    mem_c[58] = 8'b00000000;
    mem_c[59] = 8'b00000000;
    mem_c[60] = 8'b00000000;
    mem_c[61] = 8'b00000000;
    mem_c[62] = 8'b00000000;
    mem_c[63] = 8'b00000000;
    mem_c[64] = 8'b00000000;
    mem_c[65] = 8'b00000000;
    mem_c[66] = 8'b00000000;
    mem_c[67] = 8'b00000000;
    mem_c[68] = 8'b00000000;
    mem_c[69] = 8'b00000000;
    mem_c[70] = 8'b00000000;
    mem_c[71] = 8'b00000000;
    mem_c[72] = 8'b00000000;
    mem_c[73] = 8'b00000000;
    mem_c[74] = 8'b00000000;
    mem_c[75] = 8'b00000000;
    mem_c[76] = 8'b00000000;
    mem_c[77] = 8'b00000000;
    mem_c[78] = 8'b00000000;
    mem_c[79] = 8'b00000000;
    mem_c[80] = 8'b00000000;
    mem_c[81] = 8'b00000000;
    mem_c[82] = 8'b00000000;
    mem_c[83] = 8'b00000000;
    mem_c[84] = 8'b00000000;
    mem_c[85] = 8'b00000000;
    mem_c[86] = 8'b00000000;
    mem_c[87] = 8'b00000000;
    mem_c[88] = 8'b00000000;
    mem_c[89] = 8'b00000000;
    mem_c[90] = 8'b00000000;
    mem_c[91] = 8'b00000000;
    mem_c[92] = 8'b00000000;
    mem_c[93] = 8'b00111000;
    mem_c[94] = 8'b00000000;
    mem_c[95] = 8'b00000000;
    mem_c[96] = 8'b00000000;
    mem_c[97] = 8'b00000000;
    mem_c[98] = 8'b00111100;
    mem_c[99] = 8'b00000000;
    mem_c[100] = 8'b00000000;
    mem_c[101] = 8'b00000000;
    mem_c[102] = 8'b00000000;
    mem_c[103] = 8'b00000000;
    mem_c[104] = 8'b00000000;
    mem_c[105] = 8'b00000000;
    mem_c[106] = 8'b00000000;
    mem_c[107] = 8'b00000000;
    mem_c[108] = 8'b00000000;
    mem_c[109] = 8'b00111111;
    mem_c[110] = 8'b00000000;
    mem_c[111] = 8'b00000000;
    mem_c[112] = 8'b00000000;
    mem_c[113] = 8'b00000000;
    mem_c[114] = 8'b11111100;
    mem_c[115] = 8'b00000000;
    mem_c[116] = 8'b00000000;
    mem_c[117] = 8'b00000000;
    mem_c[118] = 8'b00000000;
    mem_c[119] = 8'b00000000;
    mem_c[120] = 8'b00000000;
    mem_c[121] = 8'b00000000;
    mem_c[122] = 8'b00000000;
    mem_c[123] = 8'b00000000;
    mem_c[124] = 8'b11000000;
    mem_c[125] = 8'b00111111;
    mem_c[126] = 8'b00000000;
    mem_c[127] = 8'b00000000;
    mem_c[128] = 8'b00000000;
    mem_c[129] = 8'b00000000;
    mem_c[130] = 8'b11111100;
    mem_c[131] = 8'b00000011;
    mem_c[132] = 8'b00000000;
    mem_c[133] = 8'b00000000;
    mem_c[134] = 8'b00000000;
    mem_c[135] = 8'b00000000;
    mem_c[136] = 8'b00000000;
    mem_c[137] = 8'b00000000;
    mem_c[138] = 8'b00000000;
    mem_c[139] = 8'b00000000;
    mem_c[140] = 8'b11110000;
    mem_c[141] = 8'b01111111;
    mem_c[142] = 8'b00000000;
    mem_c[143] = 8'b00000000;
    mem_c[144] = 8'b00000000;
    mem_c[145] = 8'b00000000;
    mem_c[146] = 8'b11111110;
    mem_c[147] = 8'b00000111;
    mem_c[148] = 8'b00000000;
    mem_c[149] = 8'b00000000;
    mem_c[150] = 8'b00000000;
    mem_c[151] = 8'b00000000;
    mem_c[152] = 8'b00000000;
    mem_c[153] = 8'b00000000;
    mem_c[154] = 8'b00000000;
    mem_c[155] = 8'b00000000;
    mem_c[156] = 8'b11111100;
    mem_c[157] = 8'b01111111;
    mem_c[158] = 8'b00000000;
    mem_c[159] = 8'b00000000;
    mem_c[160] = 8'b00000000;
    mem_c[161] = 8'b00000000;
    mem_c[162] = 8'b11111110;
    mem_c[163] = 8'b00001111;
    mem_c[164] = 8'b00000000;
    mem_c[165] = 8'b00000000;
    mem_c[166] = 8'b00000000;
    mem_c[167] = 8'b00000000;
    mem_c[168] = 8'b00000000;
    mem_c[169] = 8'b00000000;
    mem_c[170] = 8'b00000000;
    mem_c[171] = 8'b00000000;
    mem_c[172] = 8'b11111111;
    mem_c[173] = 8'b01111111;
    mem_c[174] = 8'b00000000;
    mem_c[175] = 8'b00000000;
    mem_c[176] = 8'b00000000;
    mem_c[177] = 8'b00000000;
    mem_c[178] = 8'b11111110;
    mem_c[179] = 8'b00111111;
    mem_c[180] = 8'b00000000;
    mem_c[181] = 8'b00000000;
    mem_c[182] = 8'b00000000;
    mem_c[183] = 8'b00000000;
    mem_c[184] = 8'b00000000;
    mem_c[185] = 8'b00000000;
    mem_c[186] = 8'b00000000;
    mem_c[187] = 8'b11000000;
    mem_c[188] = 8'b11111111;
    mem_c[189] = 8'b11111111;
    mem_c[190] = 8'b00000000;
    mem_c[191] = 8'b00000000;
    mem_c[192] = 8'b00000000;
    mem_c[193] = 8'b00000000;
    mem_c[194] = 8'b11111111;
    mem_c[195] = 8'b01111111;
    mem_c[196] = 8'b00000000;
    mem_c[197] = 8'b00000000;
    mem_c[198] = 8'b00000000;
    mem_c[199] = 8'b00000000;
    mem_c[200] = 8'b00000000;
    mem_c[201] = 8'b00000000;
    mem_c[202] = 8'b00000000;
    mem_c[203] = 8'b11100000;
    mem_c[204] = 8'b11111111;
    mem_c[205] = 8'b11111111;
    mem_c[206] = 8'b00000000;
    mem_c[207] = 8'b00000000;
    mem_c[208] = 8'b00000000;
    mem_c[209] = 8'b00000000;
    mem_c[210] = 8'b11111111;
    mem_c[211] = 8'b11111111;
    mem_c[212] = 8'b00000000;
    mem_c[213] = 8'b00000000;
    mem_c[214] = 8'b11100000;
    mem_c[215] = 8'b00000001;
    mem_c[216] = 8'b00000000;
    mem_c[217] = 8'b00000000;
    mem_c[218] = 8'b00000000;
    mem_c[219] = 8'b11110000;
    mem_c[220] = 8'b11111111;
    mem_c[221] = 8'b11111111;
    mem_c[222] = 8'b00000000;
    mem_c[223] = 8'b00000000;
    mem_c[224] = 8'b00000000;
    mem_c[225] = 8'b00000000;
    mem_c[226] = 8'b11111111;
    mem_c[227] = 8'b11111111;
    mem_c[228] = 8'b00000011;
    mem_c[229] = 8'b00000000;
    mem_c[230] = 8'b11100000;
    mem_c[231] = 8'b00011111;
    mem_c[232] = 8'b00000000;
    mem_c[233] = 8'b00000000;
    mem_c[234] = 8'b00000000;
    mem_c[235] = 8'b11111000;
    mem_c[236] = 8'b11111111;
    mem_c[237] = 8'b11111111;
    mem_c[238] = 8'b00000000;
    mem_c[239] = 8'b00000000;
    mem_c[240] = 8'b00000000;
    mem_c[241] = 8'b00000000;
    mem_c[242] = 8'b11111111;
    mem_c[243] = 8'b11111111;
    mem_c[244] = 8'b00000111;
    mem_c[245] = 8'b00000000;
    mem_c[246] = 8'b11000000;
    mem_c[247] = 8'b11111111;
    mem_c[248] = 8'b00000000;
    mem_c[249] = 8'b00000000;
    mem_c[250] = 8'b00000000;
    mem_c[251] = 8'b11111100;
    mem_c[252] = 8'b11111111;
    mem_c[253] = 8'b11111111;
    mem_c[254] = 8'b00000001;
    mem_c[255] = 8'b00000000;
    mem_c[256] = 8'b00000000;
    mem_c[257] = 8'b00000000;
    mem_c[258] = 8'b11111111;
    mem_c[259] = 8'b11111111;
    mem_c[260] = 8'b00001111;
    mem_c[261] = 8'b00000000;
    mem_c[262] = 8'b11000000;
    mem_c[263] = 8'b11111111;
    mem_c[264] = 8'b00000011;
    mem_c[265] = 8'b00000000;
    mem_c[266] = 8'b00000000;
    mem_c[267] = 8'b11111110;
    mem_c[268] = 8'b11111111;
    mem_c[269] = 8'b11111111;
    mem_c[270] = 8'b00000001;
    mem_c[271] = 8'b00000000;
    mem_c[272] = 8'b00000000;
    mem_c[273] = 8'b10000000;
    mem_c[274] = 8'b11111111;
    mem_c[275] = 8'b11111111;
    mem_c[276] = 8'b00011111;
    mem_c[277] = 8'b00000000;
    mem_c[278] = 8'b10000000;
    mem_c[279] = 8'b11111111;
    mem_c[280] = 8'b00001111;
    mem_c[281] = 8'b00000000;
    mem_c[282] = 8'b10000000;
    mem_c[283] = 8'b11111111;
    mem_c[284] = 8'b11111111;
    mem_c[285] = 8'b11111111;
    mem_c[286] = 8'b00000001;
    mem_c[287] = 8'b00000000;
    mem_c[288] = 8'b00000000;
    mem_c[289] = 8'b10000000;
    mem_c[290] = 8'b11111111;
    mem_c[291] = 8'b11111111;
    mem_c[292] = 8'b00111111;
    mem_c[293] = 8'b00000000;
    mem_c[294] = 8'b10000000;
    mem_c[295] = 8'b11111111;
    mem_c[296] = 8'b00111111;
    mem_c[297] = 8'b00000000;
    mem_c[298] = 8'b10000000;
    mem_c[299] = 8'b11111111;
    mem_c[300] = 8'b11111111;
    mem_c[301] = 8'b11111111;
    mem_c[302] = 8'b00000001;
    mem_c[303] = 8'b00000000;
    mem_c[304] = 8'b00000000;
    mem_c[305] = 8'b10000000;
    mem_c[306] = 8'b11111111;
    mem_c[307] = 8'b11111111;
    mem_c[308] = 8'b01111111;
    mem_c[309] = 8'b00000000;
    mem_c[310] = 8'b00000000;
    mem_c[311] = 8'b11111111;
    mem_c[312] = 8'b11111111;
    mem_c[313] = 8'b00000000;
    mem_c[314] = 8'b11000000;
    mem_c[315] = 8'b11111111;
    mem_c[316] = 8'b11111111;
    mem_c[317] = 8'b11111111;
    mem_c[318] = 8'b00000011;
    mem_c[319] = 8'b00000000;
    mem_c[320] = 8'b00000000;
    mem_c[321] = 8'b10000000;
    mem_c[322] = 8'b11111111;
    mem_c[323] = 8'b11111111;
    mem_c[324] = 8'b11111111;
    mem_c[325] = 8'b00000000;
    mem_c[326] = 8'b00000000;
    mem_c[327] = 8'b11111110;
    mem_c[328] = 8'b11111111;
    mem_c[329] = 8'b00000001;
    mem_c[330] = 8'b11000000;
    mem_c[331] = 8'b11111111;
    mem_c[332] = 8'b11111111;
    mem_c[333] = 8'b11111111;
    mem_c[334] = 8'b00000011;
    mem_c[335] = 8'b00000000;
    mem_c[336] = 8'b00000000;
    mem_c[337] = 8'b10000000;
    mem_c[338] = 8'b11111111;
    mem_c[339] = 8'b11111111;
    mem_c[340] = 8'b11111111;
    mem_c[341] = 8'b00000001;
    mem_c[342] = 8'b00000000;
    mem_c[343] = 8'b11111100;
    mem_c[344] = 8'b11111111;
    mem_c[345] = 8'b00000111;
    mem_c[346] = 8'b11100000;
    mem_c[347] = 8'b11111111;
    mem_c[348] = 8'b11111111;
    mem_c[349] = 8'b11111111;
    mem_c[350] = 8'b00000011;
    mem_c[351] = 8'b00000000;
    mem_c[352] = 8'b00000000;
    mem_c[353] = 8'b11000000;
    mem_c[354] = 8'b11111111;
    mem_c[355] = 8'b11111111;
    mem_c[356] = 8'b11111111;
    mem_c[357] = 8'b00000011;
    mem_c[358] = 8'b00000000;
    mem_c[359] = 8'b11111000;
    mem_c[360] = 8'b11111111;
    mem_c[361] = 8'b00001111;
    mem_c[362] = 8'b11100000;
    mem_c[363] = 8'b11111111;
    mem_c[364] = 8'b11111111;
    mem_c[365] = 8'b11111111;
    mem_c[366] = 8'b00000011;
    mem_c[367] = 8'b00000000;
    mem_c[368] = 8'b00000000;
    mem_c[369] = 8'b11000000;
    mem_c[370] = 8'b11111111;
    mem_c[371] = 8'b11111111;
    mem_c[372] = 8'b11111111;
    mem_c[373] = 8'b00000111;
    mem_c[374] = 8'b00000000;
    mem_c[375] = 8'b11111000;
    mem_c[376] = 8'b11111111;
    mem_c[377] = 8'b00011111;
    mem_c[378] = 8'b11110000;
    mem_c[379] = 8'b11111111;
    mem_c[380] = 8'b11111111;
    mem_c[381] = 8'b11111111;
    mem_c[382] = 8'b00000111;
    mem_c[383] = 8'b00000000;
    mem_c[384] = 8'b00000000;
    mem_c[385] = 8'b11000000;
    mem_c[386] = 8'b11111111;
    mem_c[387] = 8'b11111111;
    mem_c[388] = 8'b11111111;
    mem_c[389] = 8'b00001111;
    mem_c[390] = 8'b00000000;
    mem_c[391] = 8'b11110000;
    mem_c[392] = 8'b11111111;
    mem_c[393] = 8'b00111111;
    mem_c[394] = 8'b11110000;
    mem_c[395] = 8'b11111111;
    mem_c[396] = 8'b11111111;
    mem_c[397] = 8'b11111111;
    mem_c[398] = 8'b00000111;
    mem_c[399] = 8'b00000000;
    mem_c[400] = 8'b00000000;
    mem_c[401] = 8'b11000000;
    mem_c[402] = 8'b11111111;
    mem_c[403] = 8'b11111111;
    mem_c[404] = 8'b11111111;
    mem_c[405] = 8'b00001111;
    mem_c[406] = 8'b00000000;
    mem_c[407] = 8'b11110000;
    mem_c[408] = 8'b11111111;
    mem_c[409] = 8'b01111111;
    mem_c[410] = 8'b11111000;
    mem_c[411] = 8'b11111111;
    mem_c[412] = 8'b11111111;
    mem_c[413] = 8'b11111111;
    mem_c[414] = 8'b00000111;
    mem_c[415] = 8'b00000000;
    mem_c[416] = 8'b00000000;
    mem_c[417] = 8'b11000000;
    mem_c[418] = 8'b11111111;
    mem_c[419] = 8'b11111111;
    mem_c[420] = 8'b11111111;
    mem_c[421] = 8'b00011111;
    mem_c[422] = 8'b00000000;
    mem_c[423] = 8'b11110000;
    mem_c[424] = 8'b11111111;
    mem_c[425] = 8'b11111111;
    mem_c[426] = 8'b11111000;
    mem_c[427] = 8'b11111111;
    mem_c[428] = 8'b11111111;
    mem_c[429] = 8'b11111111;
    mem_c[430] = 8'b00000111;
    mem_c[431] = 8'b00000000;
    mem_c[432] = 8'b00000000;
    mem_c[433] = 8'b11000000;
    mem_c[434] = 8'b11111111;
    mem_c[435] = 8'b11111111;
    mem_c[436] = 8'b11111111;
    mem_c[437] = 8'b00111111;
    mem_c[438] = 8'b00000000;
    mem_c[439] = 8'b11111100;
    mem_c[440] = 8'b11111111;
    mem_c[441] = 8'b11111111;
    mem_c[442] = 8'b11111000;
    mem_c[443] = 8'b11111111;
    mem_c[444] = 8'b11111111;
    mem_c[445] = 8'b11111111;
    mem_c[446] = 8'b00000111;
    mem_c[447] = 8'b00000000;
    mem_c[448] = 8'b00000000;
    mem_c[449] = 8'b11000000;
    mem_c[450] = 8'b11111111;
    mem_c[451] = 8'b11111111;
    mem_c[452] = 8'b11111111;
    mem_c[453] = 8'b11111111;
    mem_c[454] = 8'b11000000;
    mem_c[455] = 8'b11111111;
    mem_c[456] = 8'b11111111;
    mem_c[457] = 8'b11111111;
    mem_c[458] = 8'b11111111;
    mem_c[459] = 8'b11111111;
    mem_c[460] = 8'b11111111;
    mem_c[461] = 8'b11111111;
    mem_c[462] = 8'b00001111;
    mem_c[463] = 8'b00000000;
    mem_c[464] = 8'b00000000;
    mem_c[465] = 8'b11000000;
    mem_c[466] = 8'b11111111;
    mem_c[467] = 8'b11111111;
    mem_c[468] = 8'b11111111;
    mem_c[469] = 8'b01111111;
    mem_c[470] = 8'b11100000;
    mem_c[471] = 8'b11111111;
    mem_c[472] = 8'b11111111;
    mem_c[473] = 8'b11111111;
    mem_c[474] = 8'b11111111;
    mem_c[475] = 8'b11111111;
    mem_c[476] = 8'b11111111;
    mem_c[477] = 8'b11111111;
    mem_c[478] = 8'b00001111;
    mem_c[479] = 8'b00000000;
    mem_c[480] = 8'b00000000;
    mem_c[481] = 8'b11100000;
    mem_c[482] = 8'b11111111;
    mem_c[483] = 8'b11111111;
    mem_c[484] = 8'b11111111;
    mem_c[485] = 8'b00111111;
    mem_c[486] = 8'b11110000;
    mem_c[487] = 8'b11111111;
    mem_c[488] = 8'b11111111;
    mem_c[489] = 8'b11111111;
    mem_c[490] = 8'b11111111;
    mem_c[491] = 8'b11111111;
    mem_c[492] = 8'b11111111;
    mem_c[493] = 8'b11111111;
    mem_c[494] = 8'b00001111;
    mem_c[495] = 8'b00000000;
    mem_c[496] = 8'b00000000;
    mem_c[497] = 8'b11100000;
    mem_c[498] = 8'b11111111;
    mem_c[499] = 8'b11111111;
    mem_c[500] = 8'b11111111;
    mem_c[501] = 8'b00011111;
    mem_c[502] = 8'b11111000;
    mem_c[503] = 8'b11111111;
    mem_c[504] = 8'b11111111;
    mem_c[505] = 8'b11111111;
    mem_c[506] = 8'b11111111;
    mem_c[507] = 8'b11111111;
    mem_c[508] = 8'b11111111;
    mem_c[509] = 8'b11111111;
    mem_c[510] = 8'b00001111;
    mem_c[511] = 8'b00000000;
    mem_c[512] = 8'b00000000;
    mem_c[513] = 8'b11100000;
    mem_c[514] = 8'b11111111;
    mem_c[515] = 8'b11111111;
    mem_c[516] = 8'b11111111;
    mem_c[517] = 8'b00011111;
    mem_c[518] = 8'b00000000;
    mem_c[519] = 8'b11000000;
    mem_c[520] = 8'b11111111;
    mem_c[521] = 8'b11111111;
    mem_c[522] = 8'b11111111;
    mem_c[523] = 8'b11111111;
    mem_c[524] = 8'b11111111;
    mem_c[525] = 8'b11111111;
    mem_c[526] = 8'b00001111;
    mem_c[527] = 8'b00000000;
    mem_c[528] = 8'b00000000;
    mem_c[529] = 8'b11100000;
    mem_c[530] = 8'b11111111;
    mem_c[531] = 8'b11111111;
    mem_c[532] = 8'b11111111;
    mem_c[533] = 8'b00011111;
    mem_c[534] = 8'b00000000;
    mem_c[535] = 8'b00000000;
    mem_c[536] = 8'b11111110;
    mem_c[537] = 8'b11111111;
    mem_c[538] = 8'b11111111;
    mem_c[539] = 8'b11111111;
    mem_c[540] = 8'b11111111;
    mem_c[541] = 8'b11111111;
    mem_c[542] = 8'b00011111;
    mem_c[543] = 8'b00000000;
    mem_c[544] = 8'b00000000;
    mem_c[545] = 8'b11100000;
    mem_c[546] = 8'b11111111;
    mem_c[547] = 8'b11111111;
    mem_c[548] = 8'b11111111;
    mem_c[549] = 8'b00011111;
    mem_c[550] = 8'b00000000;
    mem_c[551] = 8'b00000000;
    mem_c[552] = 8'b11111110;
    mem_c[553] = 8'b11111111;
    mem_c[554] = 8'b11111111;
    mem_c[555] = 8'b11111111;
    mem_c[556] = 8'b11111111;
    mem_c[557] = 8'b11111111;
    mem_c[558] = 8'b00011111;
    mem_c[559] = 8'b00000000;
    mem_c[560] = 8'b00000000;
    mem_c[561] = 8'b11100000;
    mem_c[562] = 8'b11111111;
    mem_c[563] = 8'b11111111;
    mem_c[564] = 8'b11111111;
    mem_c[565] = 8'b11111111;
    mem_c[566] = 8'b11111111;
    mem_c[567] = 8'b00000111;
    mem_c[568] = 8'b11111110;
    mem_c[569] = 8'b11111111;
    mem_c[570] = 8'b11111111;
    mem_c[571] = 8'b11111111;
    mem_c[572] = 8'b11111111;
    mem_c[573] = 8'b11111111;
    mem_c[574] = 8'b00011111;
    mem_c[575] = 8'b00000000;
    mem_c[576] = 8'b00000000;
    mem_c[577] = 8'b11100000;
    mem_c[578] = 8'b11111111;
    mem_c[579] = 8'b11111111;
    mem_c[580] = 8'b11111111;
    mem_c[581] = 8'b11111111;
    mem_c[582] = 8'b11111111;
    mem_c[583] = 8'b11111111;
    mem_c[584] = 8'b11111111;
    mem_c[585] = 8'b11111111;
    mem_c[586] = 8'b11111111;
    mem_c[587] = 8'b11111111;
    mem_c[588] = 8'b11111111;
    mem_c[589] = 8'b11111111;
    mem_c[590] = 8'b00011111;
    mem_c[591] = 8'b00000000;
    mem_c[592] = 8'b00000000;
    mem_c[593] = 8'b11110000;
    mem_c[594] = 8'b11111111;
    mem_c[595] = 8'b11111111;
    mem_c[596] = 8'b11111111;
    mem_c[597] = 8'b11111111;
    mem_c[598] = 8'b11111111;
    mem_c[599] = 8'b11111111;
    mem_c[600] = 8'b11111111;
    mem_c[601] = 8'b11111111;
    mem_c[602] = 8'b11111111;
    mem_c[603] = 8'b11111111;
    mem_c[604] = 8'b11111111;
    mem_c[605] = 8'b11111111;
    mem_c[606] = 8'b00011111;
    mem_c[607] = 8'b00000000;
    mem_c[608] = 8'b00000000;
    mem_c[609] = 8'b11110000;
    mem_c[610] = 8'b11111111;
    mem_c[611] = 8'b11111111;
    mem_c[612] = 8'b11111111;
    mem_c[613] = 8'b11111111;
    mem_c[614] = 8'b11111111;
    mem_c[615] = 8'b11111111;
    mem_c[616] = 8'b11111111;
    mem_c[617] = 8'b11111111;
    mem_c[618] = 8'b11111111;
    mem_c[619] = 8'b11111111;
    mem_c[620] = 8'b11111111;
    mem_c[621] = 8'b11111111;
    mem_c[622] = 8'b00011111;
    mem_c[623] = 8'b00000000;
    mem_c[624] = 8'b00000000;
    mem_c[625] = 8'b11110000;
    mem_c[626] = 8'b11111111;
    mem_c[627] = 8'b11111111;
    mem_c[628] = 8'b11111111;
    mem_c[629] = 8'b11111111;
    mem_c[630] = 8'b11111111;
    mem_c[631] = 8'b11111111;
    mem_c[632] = 8'b11111111;
    mem_c[633] = 8'b11111111;
    mem_c[634] = 8'b11111111;
    mem_c[635] = 8'b11111111;
    mem_c[636] = 8'b11111111;
    mem_c[637] = 8'b11111111;
    mem_c[638] = 8'b00011111;
    mem_c[639] = 8'b00000000;
    mem_c[640] = 8'b00000000;
    mem_c[641] = 8'b11100000;
    mem_c[642] = 8'b11111111;
    mem_c[643] = 8'b11111111;
    mem_c[644] = 8'b11111111;
    mem_c[645] = 8'b11111111;
    mem_c[646] = 8'b11111111;
    mem_c[647] = 8'b11111111;
    mem_c[648] = 8'b11111111;
    mem_c[649] = 8'b11111111;
    mem_c[650] = 8'b11111111;
    mem_c[651] = 8'b11111111;
    mem_c[652] = 8'b11111111;
    mem_c[653] = 8'b11111111;
    mem_c[654] = 8'b00011111;
    mem_c[655] = 8'b00000000;
    mem_c[656] = 8'b00000000;
    mem_c[657] = 8'b11100000;
    mem_c[658] = 8'b11111111;
    mem_c[659] = 8'b11111111;
    mem_c[660] = 8'b11111111;
    mem_c[661] = 8'b11111111;
    mem_c[662] = 8'b11111111;
    mem_c[663] = 8'b11111111;
    mem_c[664] = 8'b11111111;
    mem_c[665] = 8'b11111111;
    mem_c[666] = 8'b11111111;
    mem_c[667] = 8'b11111111;
    mem_c[668] = 8'b11111111;
    mem_c[669] = 8'b11111111;
    mem_c[670] = 8'b00001111;
    mem_c[671] = 8'b00000000;
    mem_c[672] = 8'b00000000;
    mem_c[673] = 8'b11100000;
    mem_c[674] = 8'b11111111;
    mem_c[675] = 8'b11111111;
    mem_c[676] = 8'b11111111;
    mem_c[677] = 8'b11111111;
    mem_c[678] = 8'b11111111;
    mem_c[679] = 8'b11111111;
    mem_c[680] = 8'b11111111;
    mem_c[681] = 8'b11111111;
    mem_c[682] = 8'b11111111;
    mem_c[683] = 8'b11111111;
    mem_c[684] = 8'b11111111;
    mem_c[685] = 8'b11111111;
    mem_c[686] = 8'b00001111;
    mem_c[687] = 8'b00000000;
    mem_c[688] = 8'b00000000;
    mem_c[689] = 8'b11100000;
    mem_c[690] = 8'b11111111;
    mem_c[691] = 8'b11111111;
    mem_c[692] = 8'b11111111;
    mem_c[693] = 8'b11111111;
    mem_c[694] = 8'b11111111;
    mem_c[695] = 8'b11111111;
    mem_c[696] = 8'b11111111;
    mem_c[697] = 8'b11111111;
    mem_c[698] = 8'b11111111;
    mem_c[699] = 8'b11111111;
    mem_c[700] = 8'b11111111;
    mem_c[701] = 8'b11111111;
    mem_c[702] = 8'b00001111;
    mem_c[703] = 8'b00000000;
    mem_c[704] = 8'b00000000;
    mem_c[705] = 8'b11000000;
    mem_c[706] = 8'b11111111;
    mem_c[707] = 8'b11111111;
    mem_c[708] = 8'b11111111;
    mem_c[709] = 8'b11111111;
    mem_c[710] = 8'b11111111;
    mem_c[711] = 8'b11111111;
    mem_c[712] = 8'b11111111;
    mem_c[713] = 8'b11111111;
    mem_c[714] = 8'b11111111;
    mem_c[715] = 8'b11111111;
    mem_c[716] = 8'b11111111;
    mem_c[717] = 8'b11111111;
    mem_c[718] = 8'b00001111;
    mem_c[719] = 8'b00000000;
    mem_c[720] = 8'b00000000;
    mem_c[721] = 8'b11000000;
    mem_c[722] = 8'b11111111;
    mem_c[723] = 8'b11111111;
    mem_c[724] = 8'b11111111;
    mem_c[725] = 8'b11111111;
    mem_c[726] = 8'b11111111;
    mem_c[727] = 8'b11111111;
    mem_c[728] = 8'b11111111;
    mem_c[729] = 8'b11111111;
    mem_c[730] = 8'b11111111;
    mem_c[731] = 8'b11111111;
    mem_c[732] = 8'b11111111;
    mem_c[733] = 8'b11111111;
    mem_c[734] = 8'b00001111;
    mem_c[735] = 8'b00000000;
    mem_c[736] = 8'b00000000;
    mem_c[737] = 8'b11000000;
    mem_c[738] = 8'b11111111;
    mem_c[739] = 8'b11111111;
    mem_c[740] = 8'b11111111;
    mem_c[741] = 8'b11111111;
    mem_c[742] = 8'b11111111;
    mem_c[743] = 8'b11111111;
    mem_c[744] = 8'b11111111;
    mem_c[745] = 8'b11111111;
    mem_c[746] = 8'b11111111;
    mem_c[747] = 8'b11111111;
    mem_c[748] = 8'b11111111;
    mem_c[749] = 8'b11111111;
    mem_c[750] = 8'b00000111;
    mem_c[751] = 8'b00000000;
    mem_c[752] = 8'b00000000;
    mem_c[753] = 8'b10000000;
    mem_c[754] = 8'b11111111;
    mem_c[755] = 8'b11111111;
    mem_c[756] = 8'b11111111;
    mem_c[757] = 8'b11111111;
    mem_c[758] = 8'b11111111;
    mem_c[759] = 8'b11111111;
    mem_c[760] = 8'b11111111;
    mem_c[761] = 8'b11111111;
    mem_c[762] = 8'b11111111;
    mem_c[763] = 8'b11111111;
    mem_c[764] = 8'b11111111;
    mem_c[765] = 8'b11111111;
    mem_c[766] = 8'b00000111;
    mem_c[767] = 8'b00000000;
    mem_c[768] = 8'b00000000;
    mem_c[769] = 8'b10000000;
    mem_c[770] = 8'b11111111;
    mem_c[771] = 8'b11111111;
    mem_c[772] = 8'b11111111;
    mem_c[773] = 8'b11111111;
    mem_c[774] = 8'b11111111;
    mem_c[775] = 8'b11111111;
    mem_c[776] = 8'b11111111;
    mem_c[777] = 8'b11111111;
    mem_c[778] = 8'b11111111;
    mem_c[779] = 8'b11111111;
    mem_c[780] = 8'b11111111;
    mem_c[781] = 8'b11111111;
    mem_c[782] = 8'b00000011;
    mem_c[783] = 8'b00000000;
    mem_c[784] = 8'b00000000;
    mem_c[785] = 8'b00000000;
    mem_c[786] = 8'b11111111;
    mem_c[787] = 8'b11111111;
    mem_c[788] = 8'b11111111;
    mem_c[789] = 8'b11111111;
    mem_c[790] = 8'b11111111;
    mem_c[791] = 8'b11111111;
    mem_c[792] = 8'b11111111;
    mem_c[793] = 8'b11111111;
    mem_c[794] = 8'b11111111;
    mem_c[795] = 8'b11111111;
    mem_c[796] = 8'b11111111;
    mem_c[797] = 8'b11111111;
    mem_c[798] = 8'b00000001;
    mem_c[799] = 8'b00000000;
    mem_c[800] = 8'b00000000;
    mem_c[801] = 8'b00000000;
    mem_c[802] = 8'b11111111;
    mem_c[803] = 8'b11111111;
    mem_c[804] = 8'b11111111;
    mem_c[805] = 8'b11111111;
    mem_c[806] = 8'b11111111;
    mem_c[807] = 8'b11111111;
    mem_c[808] = 8'b11111111;
    mem_c[809] = 8'b01111111;
    mem_c[810] = 8'b00000000;
    mem_c[811] = 8'b00000000;
    mem_c[812] = 8'b11110000;
    mem_c[813] = 8'b11111111;
    mem_c[814] = 8'b00000001;
    mem_c[815] = 8'b00000000;
    mem_c[816] = 8'b00000000;
    mem_c[817] = 8'b00000000;
    mem_c[818] = 8'b11111111;
    mem_c[819] = 8'b11111111;
    mem_c[820] = 8'b11111111;
    mem_c[821] = 8'b11111111;
    mem_c[822] = 8'b11111111;
    mem_c[823] = 8'b11111111;
    mem_c[824] = 8'b11111111;
    mem_c[825] = 8'b00011111;
    mem_c[826] = 8'b00000000;
    mem_c[827] = 8'b00000000;
    mem_c[828] = 8'b11110000;
    mem_c[829] = 8'b11111111;
    mem_c[830] = 8'b00000000;
    mem_c[831] = 8'b00000000;
    mem_c[832] = 8'b00000000;
    mem_c[833] = 8'b00000000;
    mem_c[834] = 8'b11111110;
    mem_c[835] = 8'b00000111;
    mem_c[836] = 8'b00000000;
    mem_c[837] = 8'b00000000;
    mem_c[838] = 8'b11111000;
    mem_c[839] = 8'b11111111;
    mem_c[840] = 8'b11111111;
    mem_c[841] = 8'b00000111;
    mem_c[842] = 8'b00000000;
    mem_c[843] = 8'b00000000;
    mem_c[844] = 8'b11110000;
    mem_c[845] = 8'b01111111;
    mem_c[846] = 8'b00000000;
    mem_c[847] = 8'b00000000;
    mem_c[848] = 8'b00000000;
    mem_c[849] = 8'b00000000;
    mem_c[850] = 8'b11111110;
    mem_c[851] = 8'b00000111;
    mem_c[852] = 8'b00000000;
    mem_c[853] = 8'b00000000;
    mem_c[854] = 8'b11100000;
    mem_c[855] = 8'b11111111;
    mem_c[856] = 8'b11111111;
    mem_c[857] = 8'b00000111;
    mem_c[858] = 8'b10000000;
    mem_c[859] = 8'b00001111;
    mem_c[860] = 8'b11111110;
    mem_c[861] = 8'b00111111;
    mem_c[862] = 8'b00000000;
    mem_c[863] = 8'b00000000;
    mem_c[864] = 8'b00000000;
    mem_c[865] = 8'b00000000;
    mem_c[866] = 8'b11111110;
    mem_c[867] = 8'b00000111;
    mem_c[868] = 8'b00000000;
    mem_c[869] = 8'b00000000;
    mem_c[870] = 8'b11100000;
    mem_c[871] = 8'b11111111;
    mem_c[872] = 8'b11111111;
    mem_c[873] = 8'b00000111;
    mem_c[874] = 8'b10000000;
    mem_c[875] = 8'b00001111;
    mem_c[876] = 8'b11111110;
    mem_c[877] = 8'b00011111;
    mem_c[878] = 8'b00000000;
    mem_c[879] = 8'b00000000;
    mem_c[880] = 8'b00000000;
    mem_c[881] = 8'b00000000;
    mem_c[882] = 8'b11111100;
    mem_c[883] = 8'b00111111;
    mem_c[884] = 8'b11111000;
    mem_c[885] = 8'b00000000;
    mem_c[886] = 8'b11000000;
    mem_c[887] = 8'b11111111;
    mem_c[888] = 8'b11111111;
    mem_c[889] = 8'b00000011;
    mem_c[890] = 8'b10000000;
    mem_c[891] = 8'b00011111;
    mem_c[892] = 8'b11111110;
    mem_c[893] = 8'b00001111;
    mem_c[894] = 8'b00000000;
    mem_c[895] = 8'b00000000;
    mem_c[896] = 8'b00000000;
    mem_c[897] = 8'b00000000;
    mem_c[898] = 8'b11111100;
    mem_c[899] = 8'b00011111;
    mem_c[900] = 8'b11111000;
    mem_c[901] = 8'b00000000;
    mem_c[902] = 8'b11000000;
    mem_c[903] = 8'b11111111;
    mem_c[904] = 8'b11111111;
    mem_c[905] = 8'b00000011;
    mem_c[906] = 8'b10000000;
    mem_c[907] = 8'b00111111;
    mem_c[908] = 8'b11111100;
    mem_c[909] = 8'b00001111;
    mem_c[910] = 8'b00000000;
    mem_c[911] = 8'b00000000;
    mem_c[912] = 8'b00000000;
    mem_c[913] = 8'b00000000;
    mem_c[914] = 8'b11111000;
    mem_c[915] = 8'b00011111;
    mem_c[916] = 8'b11111100;
    mem_c[917] = 8'b00000000;
    mem_c[918] = 8'b11000000;
    mem_c[919] = 8'b11111111;
    mem_c[920] = 8'b11111111;
    mem_c[921] = 8'b00000011;
    mem_c[922] = 8'b10000000;
    mem_c[923] = 8'b00111111;
    mem_c[924] = 8'b11111100;
    mem_c[925] = 8'b00000011;
    mem_c[926] = 8'b00000000;
    mem_c[927] = 8'b00000000;
    mem_c[928] = 8'b00000000;
    mem_c[929] = 8'b00000000;
    mem_c[930] = 8'b11111000;
    mem_c[931] = 8'b00001111;
    mem_c[932] = 8'b11111110;
    mem_c[933] = 8'b00000000;
    mem_c[934] = 8'b11000000;
    mem_c[935] = 8'b11111111;
    mem_c[936] = 8'b11111111;
    mem_c[937] = 8'b00000011;
    mem_c[938] = 8'b10000000;
    mem_c[939] = 8'b01111111;
    mem_c[940] = 8'b11111100;
    mem_c[941] = 8'b00000001;
    mem_c[942] = 8'b00000000;
    mem_c[943] = 8'b00000000;
    mem_c[944] = 8'b00000000;
    mem_c[945] = 8'b00000000;
    mem_c[946] = 8'b11110000;
    mem_c[947] = 8'b00001111;
    mem_c[948] = 8'b11111111;
    mem_c[949] = 8'b00000000;
    mem_c[950] = 8'b11000000;
    mem_c[951] = 8'b11111111;
    mem_c[952] = 8'b11111111;
    mem_c[953] = 8'b00000011;
    mem_c[954] = 8'b10000000;
    mem_c[955] = 8'b01111111;
    mem_c[956] = 8'b11111100;
    mem_c[957] = 8'b00000000;
    mem_c[958] = 8'b00000000;
    mem_c[959] = 8'b00000000;
    mem_c[960] = 8'b00000000;
    mem_c[961] = 8'b00000000;
    mem_c[962] = 8'b11110000;
    mem_c[963] = 8'b00001111;
    mem_c[964] = 8'b11111111;
    mem_c[965] = 8'b00000000;
    mem_c[966] = 8'b11000000;
    mem_c[967] = 8'b11111111;
    mem_c[968] = 8'b11111111;
    mem_c[969] = 8'b00000011;
    mem_c[970] = 8'b10000000;
    mem_c[971] = 8'b01111111;
    mem_c[972] = 8'b11111000;
    mem_c[973] = 8'b00000000;
    mem_c[974] = 8'b00000000;
    mem_c[975] = 8'b00000000;
    mem_c[976] = 8'b00000000;
    mem_c[977] = 8'b00000000;
    mem_c[978] = 8'b11100000;
    mem_c[979] = 8'b10000111;
    mem_c[980] = 8'b11111111;
    mem_c[981] = 8'b00000000;
    mem_c[982] = 8'b11000000;
    mem_c[983] = 8'b11111111;
    mem_c[984] = 8'b11111111;
    mem_c[985] = 8'b00000011;
    mem_c[986] = 8'b10000000;
    mem_c[987] = 8'b01111111;
    mem_c[988] = 8'b11111000;
    mem_c[989] = 8'b00000000;
    mem_c[990] = 8'b00111100;
    mem_c[991] = 8'b00000000;
    mem_c[992] = 8'b00000000;
    mem_c[993] = 8'b00000000;
    mem_c[994] = 8'b11100000;
    mem_c[995] = 8'b10000111;
    mem_c[996] = 8'b11111111;
    mem_c[997] = 8'b00000000;
    mem_c[998] = 8'b11000000;
    mem_c[999] = 8'b11111111;
    mem_c[1000] = 8'b11111111;
    mem_c[1001] = 8'b00000011;
    mem_c[1002] = 8'b10000000;
    mem_c[1003] = 8'b01111111;
    mem_c[1004] = 8'b11111000;
    mem_c[1005] = 8'b11111000;
    mem_c[1006] = 8'b00011111;
    mem_c[1007] = 8'b00000000;
    mem_c[1008] = 8'b00000000;
    mem_c[1009] = 8'b00000000;
    mem_c[1010] = 8'b00000000;
    mem_c[1011] = 8'b10000110;
    mem_c[1012] = 8'b11111111;
    mem_c[1013] = 8'b00000000;
    mem_c[1014] = 8'b11000000;
    mem_c[1015] = 8'b11111111;
    mem_c[1016] = 8'b11111111;
    mem_c[1017] = 8'b00000011;
    mem_c[1018] = 8'b10000000;
    mem_c[1019] = 8'b11111111;
    mem_c[1020] = 8'b11111000;
    mem_c[1021] = 8'b11111111;
    mem_c[1022] = 8'b00011111;
    mem_c[1023] = 8'b00000000;
    mem_c[1024] = 8'b00000000;
    mem_c[1025] = 8'b00000000;
    mem_c[1026] = 8'b00000000;
    mem_c[1027] = 8'b11000110;
    mem_c[1028] = 8'b11111111;
    mem_c[1029] = 8'b00000000;
    mem_c[1030] = 8'b11100000;
    mem_c[1031] = 8'b11111111;
    mem_c[1032] = 8'b11111111;
    mem_c[1033] = 8'b00000011;
    mem_c[1034] = 8'b10000000;
    mem_c[1035] = 8'b11111111;
    mem_c[1036] = 8'b11111000;
    mem_c[1037] = 8'b11111111;
    mem_c[1038] = 8'b00001111;
    mem_c[1039] = 8'b00000000;
    mem_c[1040] = 8'b00000000;
    mem_c[1041] = 8'b00000000;
    mem_c[1042] = 8'b00000000;
    mem_c[1043] = 8'b11000110;
    mem_c[1044] = 8'b11111111;
    mem_c[1045] = 8'b00000000;
    mem_c[1046] = 8'b11100000;
    mem_c[1047] = 8'b11111111;
    mem_c[1048] = 8'b11111111;
    mem_c[1049] = 8'b00000011;
    mem_c[1050] = 8'b10000000;
    mem_c[1051] = 8'b11111111;
    mem_c[1052] = 8'b11111000;
    mem_c[1053] = 8'b11111111;
    mem_c[1054] = 8'b00000111;
    mem_c[1055] = 8'b00000000;
    mem_c[1056] = 8'b00000000;
    mem_c[1057] = 8'b11111000;
    mem_c[1058] = 8'b11111111;
    mem_c[1059] = 8'b11000111;
    mem_c[1060] = 8'b11111111;
    mem_c[1061] = 8'b00000000;
    mem_c[1062] = 8'b11100000;
    mem_c[1063] = 8'b11111111;
    mem_c[1064] = 8'b11111111;
    mem_c[1065] = 8'b00000011;
    mem_c[1066] = 8'b10000000;
    mem_c[1067] = 8'b01111111;
    mem_c[1068] = 8'b11111000;
    mem_c[1069] = 8'b11111111;
    mem_c[1070] = 8'b00000011;
    mem_c[1071] = 8'b00000000;
    mem_c[1072] = 8'b00000000;
    mem_c[1073] = 8'b11110000;
    mem_c[1074] = 8'b11111111;
    mem_c[1075] = 8'b10000111;
    mem_c[1076] = 8'b11111111;
    mem_c[1077] = 8'b00000001;
    mem_c[1078] = 8'b11110000;
    mem_c[1079] = 8'b11111111;
    mem_c[1080] = 8'b11111111;
    mem_c[1081] = 8'b00000111;
    mem_c[1082] = 8'b11000000;
    mem_c[1083] = 8'b01111111;
    mem_c[1084] = 8'b11111000;
    mem_c[1085] = 8'b11111111;
    mem_c[1086] = 8'b00000001;
    mem_c[1087] = 8'b00000000;
    mem_c[1088] = 8'b00000000;
    mem_c[1089] = 8'b11100000;
    mem_c[1090] = 8'b11111111;
    mem_c[1091] = 8'b10000111;
    mem_c[1092] = 8'b11111111;
    mem_c[1093] = 8'b00000001;
    mem_c[1094] = 8'b11110000;
    mem_c[1095] = 8'b11111111;
    mem_c[1096] = 8'b11111111;
    mem_c[1097] = 8'b00000111;
    mem_c[1098] = 8'b11000000;
    mem_c[1099] = 8'b01111111;
    mem_c[1100] = 8'b11111000;
    mem_c[1101] = 8'b01111111;
    mem_c[1102] = 8'b00000000;
    mem_c[1103] = 8'b00000000;
    mem_c[1104] = 8'b00000000;
    mem_c[1105] = 8'b11000000;
    mem_c[1106] = 8'b11111111;
    mem_c[1107] = 8'b10000111;
    mem_c[1108] = 8'b11111111;
    mem_c[1109] = 8'b00000011;
    mem_c[1110] = 8'b11111000;
    mem_c[1111] = 8'b11111111;
    mem_c[1112] = 8'b11111111;
    mem_c[1113] = 8'b00001111;
    mem_c[1114] = 8'b11100000;
    mem_c[1115] = 8'b01111111;
    mem_c[1116] = 8'b11111100;
    mem_c[1117] = 8'b01111111;
    mem_c[1118] = 8'b00000000;
    mem_c[1119] = 8'b00000000;
    mem_c[1120] = 8'b00000000;
    mem_c[1121] = 8'b10000000;
    mem_c[1122] = 8'b11111111;
    mem_c[1123] = 8'b00001111;
    mem_c[1124] = 8'b11111111;
    mem_c[1125] = 8'b00000011;
    mem_c[1126] = 8'b11111100;
    mem_c[1127] = 8'b11111111;
    mem_c[1128] = 8'b11111111;
    mem_c[1129] = 8'b00111111;
    mem_c[1130] = 8'b11111000;
    mem_c[1131] = 8'b01111111;
    mem_c[1132] = 8'b11111100;
    mem_c[1133] = 8'b00111111;
    mem_c[1134] = 8'b00000000;
    mem_c[1135] = 8'b00000000;
    mem_c[1136] = 8'b00000000;
    mem_c[1137] = 8'b00000000;
    mem_c[1138] = 8'b11111111;
    mem_c[1139] = 8'b00001111;
    mem_c[1140] = 8'b11111111;
    mem_c[1141] = 8'b00000111;
    mem_c[1142] = 8'b11111110;
    mem_c[1143] = 8'b11111111;
    mem_c[1144] = 8'b11111111;
    mem_c[1145] = 8'b11111111;
    mem_c[1146] = 8'b11111111;
    mem_c[1147] = 8'b11111111;
    mem_c[1148] = 8'b11111111;
    mem_c[1149] = 8'b00011111;
    mem_c[1150] = 8'b00000000;
    mem_c[1151] = 8'b00000000;
    mem_c[1152] = 8'b00000000;
    mem_c[1153] = 8'b00000000;
    mem_c[1154] = 8'b11111110;
    mem_c[1155] = 8'b00001111;
    mem_c[1156] = 8'b11111111;
    mem_c[1157] = 8'b11111111;
    mem_c[1158] = 8'b11111111;
    mem_c[1159] = 8'b00000000;
    mem_c[1160] = 8'b11111111;
    mem_c[1161] = 8'b11111111;
    mem_c[1162] = 8'b11111111;
    mem_c[1163] = 8'b11111111;
    mem_c[1164] = 8'b11111111;
    mem_c[1165] = 8'b00001111;
    mem_c[1166] = 8'b00000000;
    mem_c[1167] = 8'b00000000;
    mem_c[1168] = 8'b00000000;
    mem_c[1169] = 8'b00000000;
    mem_c[1170] = 8'b11111100;
    mem_c[1171] = 8'b00011111;
    mem_c[1172] = 8'b11111111;
    mem_c[1173] = 8'b11111111;
    mem_c[1174] = 8'b11111111;
    mem_c[1175] = 8'b00000000;
    mem_c[1176] = 8'b11111111;
    mem_c[1177] = 8'b11111111;
    mem_c[1178] = 8'b11111111;
    mem_c[1179] = 8'b10000111;
    mem_c[1180] = 8'b11111111;
    mem_c[1181] = 8'b00001111;
    mem_c[1182] = 8'b00000000;
    mem_c[1183] = 8'b00000000;
    mem_c[1184] = 8'b00000000;
    mem_c[1185] = 8'b00000000;
    mem_c[1186] = 8'b11111000;
    mem_c[1187] = 8'b11110000;
    mem_c[1188] = 8'b11111111;
    mem_c[1189] = 8'b11111111;
    mem_c[1190] = 8'b11111111;
    mem_c[1191] = 8'b00000000;
    mem_c[1192] = 8'b11111111;
    mem_c[1193] = 8'b11111111;
    mem_c[1194] = 8'b11111111;
    mem_c[1195] = 8'b10000001;
    mem_c[1196] = 8'b11000011;
    mem_c[1197] = 8'b00001111;
    mem_c[1198] = 8'b00000000;
    mem_c[1199] = 8'b00000000;
    mem_c[1200] = 8'b00000000;
    mem_c[1201] = 8'b00000000;
    mem_c[1202] = 8'b01111000;
    mem_c[1203] = 8'b11100000;
    mem_c[1204] = 8'b11111111;
    mem_c[1205] = 8'b11111111;
    mem_c[1206] = 8'b11111111;
    mem_c[1207] = 8'b11111111;
    mem_c[1208] = 8'b11111111;
    mem_c[1209] = 8'b11111111;
    mem_c[1210] = 8'b11111111;
    mem_c[1211] = 8'b10000000;
    mem_c[1212] = 8'b11000001;
    mem_c[1213] = 8'b00001111;
    mem_c[1214] = 8'b00000000;
    mem_c[1215] = 8'b00000000;
    mem_c[1216] = 8'b00000000;
    mem_c[1217] = 8'b00000000;
    mem_c[1218] = 8'b00011000;
    mem_c[1219] = 8'b11100000;
    mem_c[1220] = 8'b11110001;
    mem_c[1221] = 8'b11111111;
    mem_c[1222] = 8'b11111111;
    mem_c[1223] = 8'b11111111;
    mem_c[1224] = 8'b11111111;
    mem_c[1225] = 8'b11111111;
    mem_c[1226] = 8'b01111111;
    mem_c[1227] = 8'b00000000;
    mem_c[1228] = 8'b11000000;
    mem_c[1229] = 8'b00011111;
    mem_c[1230] = 8'b00000000;
    mem_c[1231] = 8'b00000000;
    mem_c[1232] = 8'b00000000;
    mem_c[1233] = 8'b00000000;
    mem_c[1234] = 8'b00001000;
    mem_c[1235] = 8'b11000000;
    mem_c[1236] = 8'b11110000;
    mem_c[1237] = 8'b11111111;
    mem_c[1238] = 8'b11111111;
    mem_c[1239] = 8'b11111111;
    mem_c[1240] = 8'b11111111;
    mem_c[1241] = 8'b11111111;
    mem_c[1242] = 8'b00111111;
    mem_c[1243] = 8'b00000000;
    mem_c[1244] = 8'b11100000;
    mem_c[1245] = 8'b00111111;
    mem_c[1246] = 8'b00000000;
    mem_c[1247] = 8'b00000000;
    mem_c[1248] = 8'b00000000;
    mem_c[1249] = 8'b00000000;
    mem_c[1250] = 8'b00001100;
    mem_c[1251] = 8'b00000010;
    mem_c[1252] = 8'b11110000;
    mem_c[1253] = 8'b11111111;
    mem_c[1254] = 8'b11111111;
    mem_c[1255] = 8'b11111111;
    mem_c[1256] = 8'b11111111;
    mem_c[1257] = 8'b11111111;
    mem_c[1258] = 8'b00111111;
    mem_c[1259] = 8'b00001000;
    mem_c[1260] = 8'b11110000;
    mem_c[1261] = 8'b01111111;
    mem_c[1262] = 8'b00000000;
    mem_c[1263] = 8'b00000000;
    mem_c[1264] = 8'b00000000;
    mem_c[1265] = 8'b00000000;
    mem_c[1266] = 8'b00001100;
    mem_c[1267] = 8'b00000011;
    mem_c[1268] = 8'b11110000;
    mem_c[1269] = 8'b11111111;
    mem_c[1270] = 8'b11111111;
    mem_c[1271] = 8'b11111111;
    mem_c[1272] = 8'b11111111;
    mem_c[1273] = 8'b11100011;
    mem_c[1274] = 8'b00111111;
    mem_c[1275] = 8'b00001100;
    mem_c[1276] = 8'b11111100;
    mem_c[1277] = 8'b11111111;
    mem_c[1278] = 8'b00000000;
    mem_c[1279] = 8'b00000000;
    mem_c[1280] = 8'b00000000;
    mem_c[1281] = 8'b00000000;
    mem_c[1282] = 8'b11111110;
    mem_c[1283] = 8'b00000111;
    mem_c[1284] = 8'b11111000;
    mem_c[1285] = 8'b11111111;
    mem_c[1286] = 8'b11111111;
    mem_c[1287] = 8'b00011111;
    mem_c[1288] = 8'b11111111;
    mem_c[1289] = 8'b11100000;
    mem_c[1290] = 8'b11111111;
    mem_c[1291] = 8'b00001111;
    mem_c[1292] = 8'b11111110;
    mem_c[1293] = 8'b11111111;
    mem_c[1294] = 8'b00000001;
    mem_c[1295] = 8'b00000000;
    mem_c[1296] = 8'b00000000;
    mem_c[1297] = 8'b00000000;
    mem_c[1298] = 8'b11111110;
    mem_c[1299] = 8'b00000111;
    mem_c[1300] = 8'b11111110;
    mem_c[1301] = 8'b11111111;
    mem_c[1302] = 8'b11111111;
    mem_c[1303] = 8'b00001111;
    mem_c[1304] = 8'b01111110;
    mem_c[1305] = 8'b11100000;
    mem_c[1306] = 8'b11111111;
    mem_c[1307] = 8'b00001111;
    mem_c[1308] = 8'b11111111;
    mem_c[1309] = 8'b11111111;
    mem_c[1310] = 8'b00000001;
    mem_c[1311] = 8'b00000000;
    mem_c[1312] = 8'b00000000;
    mem_c[1313] = 8'b00000000;
    mem_c[1314] = 8'b11111111;
    mem_c[1315] = 8'b11111111;
    mem_c[1316] = 8'b11111111;
    mem_c[1317] = 8'b11111111;
    mem_c[1318] = 8'b11111111;
    mem_c[1319] = 8'b00000111;
    mem_c[1320] = 8'b00000000;
    mem_c[1321] = 8'b11100000;
    mem_c[1322] = 8'b11111111;
    mem_c[1323] = 8'b11111111;
    mem_c[1324] = 8'b11111111;
    mem_c[1325] = 8'b11111111;
    mem_c[1326] = 8'b00000011;
    mem_c[1327] = 8'b00000000;
    mem_c[1328] = 8'b00000000;
    mem_c[1329] = 8'b00000000;
    mem_c[1330] = 8'b11111111;
    mem_c[1331] = 8'b11111111;
    mem_c[1332] = 8'b11111111;
    mem_c[1333] = 8'b11111111;
    mem_c[1334] = 8'b10000011;
    mem_c[1335] = 8'b00000001;
    mem_c[1336] = 8'b00000000;
    mem_c[1337] = 8'b11111000;
    mem_c[1338] = 8'b11111111;
    mem_c[1339] = 8'b11111111;
    mem_c[1340] = 8'b11111111;
    mem_c[1341] = 8'b11111111;
    mem_c[1342] = 8'b00000011;
    mem_c[1343] = 8'b00000000;
    mem_c[1344] = 8'b00000000;
    mem_c[1345] = 8'b10000000;
    mem_c[1346] = 8'b11111111;
    mem_c[1347] = 8'b11111111;
    mem_c[1348] = 8'b11111111;
    mem_c[1349] = 8'b11111111;
    mem_c[1350] = 8'b00000011;
    mem_c[1351] = 8'b00000000;
    mem_c[1352] = 8'b00000000;
    mem_c[1353] = 8'b11111100;
    mem_c[1354] = 8'b11111111;
    mem_c[1355] = 8'b11111111;
    mem_c[1356] = 8'b11111111;
    mem_c[1357] = 8'b11111111;
    mem_c[1358] = 8'b00000000;
    mem_c[1359] = 8'b00000000;
    mem_c[1360] = 8'b00000000;
    mem_c[1361] = 8'b10000000;
    mem_c[1362] = 8'b11111111;
    mem_c[1363] = 8'b11111111;
    mem_c[1364] = 8'b11111111;
    mem_c[1365] = 8'b11111111;
    mem_c[1366] = 8'b00000011;
    mem_c[1367] = 8'b11000000;
    mem_c[1368] = 8'b10000001;
    mem_c[1369] = 8'b11111111;
    mem_c[1370] = 8'b11111111;
    mem_c[1371] = 8'b11111111;
    mem_c[1372] = 8'b11110000;
    mem_c[1373] = 8'b00111111;
    mem_c[1374] = 8'b00000000;
    mem_c[1375] = 8'b00000000;
    mem_c[1376] = 8'b00000000;
    mem_c[1377] = 8'b10000000;
    mem_c[1378] = 8'b11111111;
    mem_c[1379] = 8'b11111111;
    mem_c[1380] = 8'b11111111;
    mem_c[1381] = 8'b11111111;
    mem_c[1382] = 8'b00001111;
    mem_c[1383] = 8'b11110000;
    mem_c[1384] = 8'b11111111;
    mem_c[1385] = 8'b11111111;
    mem_c[1386] = 8'b11111111;
    mem_c[1387] = 8'b01111111;
    mem_c[1388] = 8'b11110000;
    mem_c[1389] = 8'b00000000;
    mem_c[1390] = 8'b00000000;
    mem_c[1391] = 8'b00000000;
    mem_c[1392] = 8'b00000000;
    mem_c[1393] = 8'b00000000;
    mem_c[1394] = 8'b01111100;
    mem_c[1395] = 8'b10000000;
    mem_c[1396] = 8'b11111111;
    mem_c[1397] = 8'b11111111;
    mem_c[1398] = 8'b11111111;
    mem_c[1399] = 8'b11111111;
    mem_c[1400] = 8'b11111111;
    mem_c[1401] = 8'b11111111;
    mem_c[1402] = 8'b11111111;
    mem_c[1403] = 8'b00111111;
    mem_c[1404] = 8'b00000000;
    mem_c[1405] = 8'b00000000;
    mem_c[1406] = 8'b00000000;
    mem_c[1407] = 8'b00000000;
    mem_c[1408] = 8'b00000000;
    mem_c[1409] = 8'b00000000;
    mem_c[1410] = 8'b00000000;
    mem_c[1411] = 8'b00000000;
    mem_c[1412] = 8'b11111110;
    mem_c[1413] = 8'b11111111;
    mem_c[1414] = 8'b11111111;
    mem_c[1415] = 8'b11111111;
    mem_c[1416] = 8'b11111111;
    mem_c[1417] = 8'b11111111;
    mem_c[1418] = 8'b11111111;
    mem_c[1419] = 8'b00001111;
    mem_c[1420] = 8'b00000000;
    mem_c[1421] = 8'b00000000;
    mem_c[1422] = 8'b00000000;
    mem_c[1423] = 8'b00000000;
    mem_c[1424] = 8'b00000000;
    mem_c[1425] = 8'b00000000;
    mem_c[1426] = 8'b00000000;
    mem_c[1427] = 8'b00000000;
    mem_c[1428] = 8'b11111100;
    mem_c[1429] = 8'b11111111;
    mem_c[1430] = 8'b11111111;
    mem_c[1431] = 8'b11111111;
    mem_c[1432] = 8'b11111111;
    mem_c[1433] = 8'b11111111;
    mem_c[1434] = 8'b11111111;
    mem_c[1435] = 8'b00000011;
    mem_c[1436] = 8'b00000000;
    mem_c[1437] = 8'b00000000;
    mem_c[1438] = 8'b00000000;
    mem_c[1439] = 8'b00000000;
    mem_c[1440] = 8'b00000000;
    mem_c[1441] = 8'b00000000;
    mem_c[1442] = 8'b00000000;
    mem_c[1443] = 8'b00000000;
    mem_c[1444] = 8'b11110000;
    mem_c[1445] = 8'b11111111;
    mem_c[1446] = 8'b11111111;
    mem_c[1447] = 8'b11111111;
    mem_c[1448] = 8'b11111111;
    mem_c[1449] = 8'b11111111;
    mem_c[1450] = 8'b11111111;
    mem_c[1451] = 8'b00000000;
    mem_c[1452] = 8'b00000000;
    mem_c[1453] = 8'b00000000;
    mem_c[1454] = 8'b00000000;
    mem_c[1455] = 8'b00000000;
    mem_c[1456] = 8'b00000000;
    mem_c[1457] = 8'b00000000;
    mem_c[1458] = 8'b00000000;
    mem_c[1459] = 8'b00000000;
    mem_c[1460] = 8'b11000000;
    mem_c[1461] = 8'b11111111;
    mem_c[1462] = 8'b11111111;
    mem_c[1463] = 8'b11111111;
    mem_c[1464] = 8'b11111111;
    mem_c[1465] = 8'b11111111;
    mem_c[1466] = 8'b00011111;
    mem_c[1467] = 8'b00000000;
    mem_c[1468] = 8'b00000000;
    mem_c[1469] = 8'b00000000;
    mem_c[1470] = 8'b00000000;
    mem_c[1471] = 8'b00000000;
    mem_c[1472] = 8'b00000000;
    mem_c[1473] = 8'b00000000;
    mem_c[1474] = 8'b00000000;
    mem_c[1475] = 8'b00000000;
    mem_c[1476] = 8'b00000000;
    mem_c[1477] = 8'b11000000;
    mem_c[1478] = 8'b11111111;
    mem_c[1479] = 8'b11111111;
    mem_c[1480] = 8'b11111111;
    mem_c[1481] = 8'b11111111;
    mem_c[1482] = 8'b00000011;
    mem_c[1483] = 8'b00000000;
    mem_c[1484] = 8'b00000000;
    mem_c[1485] = 8'b00000000;
    mem_c[1486] = 8'b00000000;
    mem_c[1487] = 8'b00000000;
    mem_c[1488] = 8'b00000000;
    mem_c[1489] = 8'b00000000;
    mem_c[1490] = 8'b00000000;
    mem_c[1491] = 8'b00000000;
    mem_c[1492] = 8'b00000000;
    mem_c[1493] = 8'b00000000;
    mem_c[1494] = 8'b11111111;
    mem_c[1495] = 8'b11111111;
    mem_c[1496] = 8'b11111111;
    mem_c[1497] = 8'b11111111;
    mem_c[1498] = 8'b00000011;
    mem_c[1499] = 8'b00000000;
    mem_c[1500] = 8'b00000000;
    mem_c[1501] = 8'b00000000;
    mem_c[1502] = 8'b00000000;
    mem_c[1503] = 8'b00000000;
    mem_c[1504] = 8'b00000000;
    mem_c[1505] = 8'b00000000;
    mem_c[1506] = 8'b00000000;
    mem_c[1507] = 8'b00000000;
    mem_c[1508] = 8'b00000000;
    mem_c[1509] = 8'b00000000;
    mem_c[1510] = 8'b11000000;
    mem_c[1511] = 8'b11111111;
    mem_c[1512] = 8'b11111111;
    mem_c[1513] = 8'b11111111;
    mem_c[1514] = 8'b10000011;
    mem_c[1515] = 8'b00000001;
    mem_c[1516] = 8'b00000000;
    mem_c[1517] = 8'b00000000;
    mem_c[1518] = 8'b00000000;
    mem_c[1519] = 8'b00000000;
    mem_c[1520] = 8'b00000000;
    mem_c[1521] = 8'b00000000;
    mem_c[1522] = 8'b00000000;
    mem_c[1523] = 8'b00000000;
    mem_c[1524] = 8'b00000000;
    mem_c[1525] = 8'b00000110;
    mem_c[1526] = 8'b11000000;
    mem_c[1527] = 8'b11111111;
    mem_c[1528] = 8'b11111111;
    mem_c[1529] = 8'b11111111;
    mem_c[1530] = 8'b11111111;
    mem_c[1531] = 8'b00000001;
    mem_c[1532] = 8'b00000000;
    mem_c[1533] = 8'b00000000;
    mem_c[1534] = 8'b00000000;
    mem_c[1535] = 8'b00000000;
    mem_c[1536] = 8'b00000000;
    mem_c[1537] = 8'b00000000;
    mem_c[1538] = 8'b00000000;
    mem_c[1539] = 8'b00000000;
    mem_c[1540] = 8'b00000000;
    mem_c[1541] = 8'b00111100;
    mem_c[1542] = 8'b11000000;
    mem_c[1543] = 8'b11111111;
    mem_c[1544] = 8'b11111111;
    mem_c[1545] = 8'b11111111;
    mem_c[1546] = 8'b00111111;
    mem_c[1547] = 8'b00000000;
    mem_c[1548] = 8'b00000000;
    mem_c[1549] = 8'b00000000;
    mem_c[1550] = 8'b00000000;
    mem_c[1551] = 8'b00000000;
    mem_c[1552] = 8'b00000000;
    mem_c[1553] = 8'b00000000;
    mem_c[1554] = 8'b00000000;
    mem_c[1555] = 8'b00000000;
    mem_c[1556] = 8'b00000000;
    mem_c[1557] = 8'b11111100;
    mem_c[1558] = 8'b11111111;
    mem_c[1559] = 8'b11111111;
    mem_c[1560] = 8'b11111111;
    mem_c[1561] = 8'b11111111;
    mem_c[1562] = 8'b00111111;
    mem_c[1563] = 8'b00000000;
    mem_c[1564] = 8'b00000000;
    mem_c[1565] = 8'b00000000;
    mem_c[1566] = 8'b00000000;
    mem_c[1567] = 8'b00000000;
    mem_c[1568] = 8'b00000000;
    mem_c[1569] = 8'b00000000;
    mem_c[1570] = 8'b00000000;
    mem_c[1571] = 8'b00000000;
    mem_c[1572] = 8'b00000000;
    mem_c[1573] = 8'b11111000;
    mem_c[1574] = 8'b11111111;
    mem_c[1575] = 8'b11111111;
    mem_c[1576] = 8'b11111111;
    mem_c[1577] = 8'b11111111;
    mem_c[1578] = 8'b00111111;
    mem_c[1579] = 8'b00000000;
    mem_c[1580] = 8'b00000000;
    mem_c[1581] = 8'b00000000;
    mem_c[1582] = 8'b00000000;
    mem_c[1583] = 8'b00000000;
    mem_c[1584] = 8'b00000000;
    mem_c[1585] = 8'b00000000;
    mem_c[1586] = 8'b00000000;
    mem_c[1587] = 8'b00000000;
    mem_c[1588] = 8'b00000000;
    mem_c[1589] = 8'b11110000;
    mem_c[1590] = 8'b11111111;
    mem_c[1591] = 8'b11111111;
    mem_c[1592] = 8'b11111111;
    mem_c[1593] = 8'b11111111;
    mem_c[1594] = 8'b01111111;
    mem_c[1595] = 8'b00000000;
    mem_c[1596] = 8'b00000000;
    mem_c[1597] = 8'b00000000;
    mem_c[1598] = 8'b00000000;
    mem_c[1599] = 8'b00000000;
    mem_c[1600] = 8'b00000000;
    mem_c[1601] = 8'b00000000;
    mem_c[1602] = 8'b00000000;
    mem_c[1603] = 8'b00000000;
    mem_c[1604] = 8'b00000000;
    mem_c[1605] = 8'b11100000;
    mem_c[1606] = 8'b11111111;
    mem_c[1607] = 8'b11111111;
    mem_c[1608] = 8'b11111111;
    mem_c[1609] = 8'b11111111;
    mem_c[1610] = 8'b01111111;
    mem_c[1611] = 8'b00000000;
    mem_c[1612] = 8'b00000000;
    mem_c[1613] = 8'b00000000;
    mem_c[1614] = 8'b00000000;
    mem_c[1615] = 8'b00000000;
    mem_c[1616] = 8'b00000000;
    mem_c[1617] = 8'b00000000;
    mem_c[1618] = 8'b00000000;
    mem_c[1619] = 8'b00000000;
    mem_c[1620] = 8'b00000000;
    mem_c[1621] = 8'b11000000;
    mem_c[1622] = 8'b11111111;
    mem_c[1623] = 8'b11111111;
    mem_c[1624] = 8'b11111111;
    mem_c[1625] = 8'b11111111;
    mem_c[1626] = 8'b11111111;
    mem_c[1627] = 8'b00000000;
    mem_c[1628] = 8'b00000000;
    mem_c[1629] = 8'b00000000;
    mem_c[1630] = 8'b00000000;
    mem_c[1631] = 8'b00000000;
    mem_c[1632] = 8'b00000000;
    mem_c[1633] = 8'b00000000;
    mem_c[1634] = 8'b00000000;
    mem_c[1635] = 8'b00000000;
    mem_c[1636] = 8'b00000000;
    mem_c[1637] = 8'b10000000;
    mem_c[1638] = 8'b11111111;
    mem_c[1639] = 8'b11111111;
    mem_c[1640] = 8'b11111111;
    mem_c[1641] = 8'b11111111;
    mem_c[1642] = 8'b11111111;
    mem_c[1643] = 8'b00000001;
    mem_c[1644] = 8'b00000000;
    mem_c[1645] = 8'b00000000;
    mem_c[1646] = 8'b00000000;
    mem_c[1647] = 8'b00000000;
    mem_c[1648] = 8'b00000000;
    mem_c[1649] = 8'b00000000;
    mem_c[1650] = 8'b00000000;
    mem_c[1651] = 8'b00000000;
    mem_c[1652] = 8'b00000000;
    mem_c[1653] = 8'b10000000;
    mem_c[1654] = 8'b11111111;
    mem_c[1655] = 8'b11111111;
    mem_c[1656] = 8'b11111111;
    mem_c[1657] = 8'b11111111;
    mem_c[1658] = 8'b11111111;
    mem_c[1659] = 8'b00000001;
    mem_c[1660] = 8'b00000000;
    mem_c[1661] = 8'b00000000;
    mem_c[1662] = 8'b00000000;
    mem_c[1663] = 8'b00000000;
    mem_c[1664] = 8'b00000000;
    mem_c[1665] = 8'b00000000;
    mem_c[1666] = 8'b00000000;
    mem_c[1667] = 8'b00000000;
    mem_c[1668] = 8'b00000000;
    mem_c[1669] = 8'b10000000;
    mem_c[1670] = 8'b11111111;
    mem_c[1671] = 8'b11111111;
    mem_c[1672] = 8'b11111111;
    mem_c[1673] = 8'b11111111;
    mem_c[1674] = 8'b11111111;
    mem_c[1675] = 8'b00000011;
    mem_c[1676] = 8'b00000000;
    mem_c[1677] = 8'b00000000;
    mem_c[1678] = 8'b00000000;
    mem_c[1679] = 8'b00000000;
    mem_c[1680] = 8'b00000000;
    mem_c[1681] = 8'b00000000;
    mem_c[1682] = 8'b00000000;
    mem_c[1683] = 8'b00000000;
    mem_c[1684] = 8'b00000000;
    mem_c[1685] = 8'b10000000;
    mem_c[1686] = 8'b11111111;
    mem_c[1687] = 8'b11111111;
    mem_c[1688] = 8'b11111111;
    mem_c[1689] = 8'b11111111;
    mem_c[1690] = 8'b11111111;
    mem_c[1691] = 8'b00000011;
    mem_c[1692] = 8'b00000000;
    mem_c[1693] = 8'b00000000;
    mem_c[1694] = 8'b00000000;
    mem_c[1695] = 8'b00000000;
    mem_c[1696] = 8'b00000000;
    mem_c[1697] = 8'b00000000;
    mem_c[1698] = 8'b00000000;
    mem_c[1699] = 8'b00000000;
    mem_c[1700] = 8'b00000000;
    mem_c[1701] = 8'b10000000;
    mem_c[1702] = 8'b11111111;
    mem_c[1703] = 8'b11111111;
    mem_c[1704] = 8'b11111111;
    mem_c[1705] = 8'b11111111;
    mem_c[1706] = 8'b11111111;
    mem_c[1707] = 8'b00000011;
    mem_c[1708] = 8'b00000000;
    mem_c[1709] = 8'b00000000;
    mem_c[1710] = 8'b00000000;
    mem_c[1711] = 8'b00000000;
    mem_c[1712] = 8'b00000000;
    mem_c[1713] = 8'b00000000;
    mem_c[1714] = 8'b00000000;
    mem_c[1715] = 8'b00000000;
    mem_c[1716] = 8'b00000000;
    mem_c[1717] = 8'b11000000;
    mem_c[1718] = 8'b11111111;
    mem_c[1719] = 8'b11111111;
    mem_c[1720] = 8'b11111111;
    mem_c[1721] = 8'b11111111;
    mem_c[1722] = 8'b11111111;
    mem_c[1723] = 8'b00000111;
    mem_c[1724] = 8'b00000000;
    mem_c[1725] = 8'b00000000;
    mem_c[1726] = 8'b00000000;
    mem_c[1727] = 8'b00000000;
    mem_c[1728] = 8'b00000000;
    mem_c[1729] = 8'b00000000;
    mem_c[1730] = 8'b00000000;
    mem_c[1731] = 8'b00000000;
    mem_c[1732] = 8'b00000000;
    mem_c[1733] = 8'b11100000;
    mem_c[1734] = 8'b11111111;
    mem_c[1735] = 8'b11111111;
    mem_c[1736] = 8'b11111111;
    mem_c[1737] = 8'b11111111;
    mem_c[1738] = 8'b11111111;
    mem_c[1739] = 8'b00000111;
    mem_c[1740] = 8'b00000000;
    mem_c[1741] = 8'b00000000;
    mem_c[1742] = 8'b00000000;
    mem_c[1743] = 8'b00000000;
    mem_c[1744] = 8'b00000000;
    mem_c[1745] = 8'b00000000;
    mem_c[1746] = 8'b00000000;
    mem_c[1747] = 8'b00000000;
    mem_c[1748] = 8'b00000000;
    mem_c[1749] = 8'b11110000;
    mem_c[1750] = 8'b11111111;
    mem_c[1751] = 8'b11111111;
    mem_c[1752] = 8'b11111111;
    mem_c[1753] = 8'b11111111;
    mem_c[1754] = 8'b11111111;
    mem_c[1755] = 8'b00000111;
    mem_c[1756] = 8'b00000000;
    mem_c[1757] = 8'b00000000;
    mem_c[1758] = 8'b00000000;
    mem_c[1759] = 8'b00000000;
    mem_c[1760] = 8'b00000000;
    mem_c[1761] = 8'b00000000;
    mem_c[1762] = 8'b00000000;
    mem_c[1763] = 8'b00000000;
    mem_c[1764] = 8'b00000000;
    mem_c[1765] = 8'b11110000;
    mem_c[1766] = 8'b11111111;
    mem_c[1767] = 8'b11111111;
    mem_c[1768] = 8'b11111111;
    mem_c[1769] = 8'b11111111;
    mem_c[1770] = 8'b11111111;
    mem_c[1771] = 8'b00000111;
    mem_c[1772] = 8'b00000000;
    mem_c[1773] = 8'b00000000;
    mem_c[1774] = 8'b00000000;
    mem_c[1775] = 8'b00000000;
    mem_c[1776] = 8'b00000000;
    mem_c[1777] = 8'b00000000;
    mem_c[1778] = 8'b00000000;
    mem_c[1779] = 8'b00000000;
    mem_c[1780] = 8'b00000000;
    mem_c[1781] = 8'b00000000;
    mem_c[1782] = 8'b11111110;
    mem_c[1783] = 8'b11111111;
    mem_c[1784] = 8'b11111111;
    mem_c[1785] = 8'b11111111;
    mem_c[1786] = 8'b11111111;
    mem_c[1787] = 8'b00001111;
    mem_c[1788] = 8'b00000000;
    mem_c[1789] = 8'b00000000;
    mem_c[1790] = 8'b00000000;
    mem_c[1791] = 8'b00000000;
    mem_c[1792] = 8'b00000000;
    mem_c[1793] = 8'b00000000;
    mem_c[1794] = 8'b00000000;
    mem_c[1795] = 8'b00000000;
    mem_c[1796] = 8'b00000000;
    mem_c[1797] = 8'b00000000;
    mem_c[1798] = 8'b11111100;
    mem_c[1799] = 8'b11111111;
    mem_c[1800] = 8'b11111111;
    mem_c[1801] = 8'b11111111;
    mem_c[1802] = 8'b11111111;
    mem_c[1803] = 8'b00001111;
    mem_c[1804] = 8'b00000000;
    mem_c[1805] = 8'b00000000;
    mem_c[1806] = 8'b00000000;
    mem_c[1807] = 8'b00000000;
    mem_c[1808] = 8'b00000000;
    mem_c[1809] = 8'b00000000;
    mem_c[1810] = 8'b00000000;
    mem_c[1811] = 8'b00000000;
    mem_c[1812] = 8'b00000000;
    mem_c[1813] = 8'b00000000;
    mem_c[1814] = 8'b11111100;
    mem_c[1815] = 8'b11111111;
    mem_c[1816] = 8'b11111111;
    mem_c[1817] = 8'b11111111;
    mem_c[1818] = 8'b11111111;
    mem_c[1819] = 8'b00001111;
    mem_c[1820] = 8'b00000000;
    mem_c[1821] = 8'b00000000;
    mem_c[1822] = 8'b00000000;
    mem_c[1823] = 8'b00000000;
    mem_c[1824] = 8'b00000000;
    mem_c[1825] = 8'b00000000;
    mem_c[1826] = 8'b00000000;
    mem_c[1827] = 8'b00000000;
    mem_c[1828] = 8'b00000000;
    mem_c[1829] = 8'b00000000;
    mem_c[1830] = 8'b11111100;
    mem_c[1831] = 8'b11111111;
    mem_c[1832] = 8'b11111111;
    mem_c[1833] = 8'b11111111;
    mem_c[1834] = 8'b11111111;
    mem_c[1835] = 8'b00011111;
    mem_c[1836] = 8'b00000000;
    mem_c[1837] = 8'b00000000;
    mem_c[1838] = 8'b00000000;
    mem_c[1839] = 8'b00000000;
    mem_c[1840] = 8'b00000000;
    mem_c[1841] = 8'b00000000;
    mem_c[1842] = 8'b00000000;
    mem_c[1843] = 8'b00000000;
    mem_c[1844] = 8'b00000000;
    mem_c[1845] = 8'b00000000;
    mem_c[1846] = 8'b11111110;
    mem_c[1847] = 8'b11111111;
    mem_c[1848] = 8'b11111111;
    mem_c[1849] = 8'b11111111;
    mem_c[1850] = 8'b11111111;
    mem_c[1851] = 8'b00011111;
    mem_c[1852] = 8'b00000000;
    mem_c[1853] = 8'b00000000;
    mem_c[1854] = 8'b00000000;
    mem_c[1855] = 8'b00000000;
    mem_c[1856] = 8'b00000000;
    mem_c[1857] = 8'b00000000;
    mem_c[1858] = 8'b00000000;
    mem_c[1859] = 8'b00000000;
    mem_c[1860] = 8'b00000000;
    mem_c[1861] = 8'b00000000;
    mem_c[1862] = 8'b11111110;
    mem_c[1863] = 8'b11111111;
    mem_c[1864] = 8'b11111111;
    mem_c[1865] = 8'b11111111;
    mem_c[1866] = 8'b11111111;
    mem_c[1867] = 8'b00011111;
    mem_c[1868] = 8'b00000000;
    mem_c[1869] = 8'b00000000;
    mem_c[1870] = 8'b00000000;
    mem_c[1871] = 8'b00000000;
    mem_c[1872] = 8'b00000000;
    mem_c[1873] = 8'b00000000;
    mem_c[1874] = 8'b00000000;
    mem_c[1875] = 8'b00000000;
    mem_c[1876] = 8'b00000000;
    mem_c[1877] = 8'b00000000;
    mem_c[1878] = 8'b11111111;
    mem_c[1879] = 8'b11111111;
    mem_c[1880] = 8'b11111111;
    mem_c[1881] = 8'b11111111;
    mem_c[1882] = 8'b11111111;
    mem_c[1883] = 8'b00111111;
    mem_c[1884] = 8'b00000000;
    mem_c[1885] = 8'b00000000;
    mem_c[1886] = 8'b00000000;
    mem_c[1887] = 8'b00000000;
    mem_c[1888] = 8'b00000000;
    mem_c[1889] = 8'b00000000;
    mem_c[1890] = 8'b00000000;
    mem_c[1891] = 8'b00000000;
    mem_c[1892] = 8'b00000000;
    mem_c[1893] = 8'b00000000;
    mem_c[1894] = 8'b11111111;
    mem_c[1895] = 8'b11111111;
    mem_c[1896] = 8'b11111111;
    mem_c[1897] = 8'b11111111;
    mem_c[1898] = 8'b11111111;
    mem_c[1899] = 8'b00111111;
    mem_c[1900] = 8'b00000000;
    mem_c[1901] = 8'b00000000;
    mem_c[1902] = 8'b00000000;
    mem_c[1903] = 8'b00000000;
    mem_c[1904] = 8'b00000000;
    mem_c[1905] = 8'b00000000;
    mem_c[1906] = 8'b00000000;
    mem_c[1907] = 8'b00000000;
    mem_c[1908] = 8'b00000000;
    mem_c[1909] = 8'b10000000;
    mem_c[1910] = 8'b11111111;
    mem_c[1911] = 8'b11111111;
    mem_c[1912] = 8'b11111111;
    mem_c[1913] = 8'b11111111;
    mem_c[1914] = 8'b11111111;
    mem_c[1915] = 8'b00111111;
    mem_c[1916] = 8'b00000000;
    mem_c[1917] = 8'b00000000;
    mem_c[1918] = 8'b00000000;
    mem_c[1919] = 8'b00000000;
    mem_c[1920] = 8'b00000000;
    mem_c[1921] = 8'b00000000;
    mem_c[1922] = 8'b00000000;
    mem_c[1923] = 8'b00000000;
    mem_c[1924] = 8'b00000000;
    mem_c[1925] = 8'b10000000;
    mem_c[1926] = 8'b11111111;
    mem_c[1927] = 8'b11111111;
    mem_c[1928] = 8'b11111111;
    mem_c[1929] = 8'b11111111;
    mem_c[1930] = 8'b11111111;
    mem_c[1931] = 8'b00111111;
    mem_c[1932] = 8'b00000000;
    mem_c[1933] = 8'b00000000;
    mem_c[1934] = 8'b00000000;
    mem_c[1935] = 8'b00000000;
    mem_c[1936] = 8'b00000000;
    mem_c[1937] = 8'b00000000;
    mem_c[1938] = 8'b00000000;
    mem_c[1939] = 8'b00000000;
    mem_c[1940] = 8'b00000000;
    mem_c[1941] = 8'b10000000;
    mem_c[1942] = 8'b11111111;
    mem_c[1943] = 8'b11111111;
    mem_c[1944] = 8'b11111111;
    mem_c[1945] = 8'b11111111;
    mem_c[1946] = 8'b11111111;
    mem_c[1947] = 8'b00111111;
    mem_c[1948] = 8'b00000000;
    mem_c[1949] = 8'b00000000;
    mem_c[1950] = 8'b00000000;
    mem_c[1951] = 8'b00000000;
    mem_c[1952] = 8'b00000000;
    mem_c[1953] = 8'b00000000;
    mem_c[1954] = 8'b00000000;
    mem_c[1955] = 8'b00000000;
    mem_c[1956] = 8'b00000000;
    mem_c[1957] = 8'b11000000;
    mem_c[1958] = 8'b11111111;
    mem_c[1959] = 8'b11111111;
    mem_c[1960] = 8'b11111111;
    mem_c[1961] = 8'b11111111;
    mem_c[1962] = 8'b11111111;
    mem_c[1963] = 8'b01111111;
    mem_c[1964] = 8'b00000000;
    mem_c[1965] = 8'b00000000;
    mem_c[1966] = 8'b00000000;
    mem_c[1967] = 8'b00000000;
    mem_c[1968] = 8'b00000000;
    mem_c[1969] = 8'b00000000;
    mem_c[1970] = 8'b00000000;
    mem_c[1971] = 8'b00000000;
    mem_c[1972] = 8'b00000000;
    mem_c[1973] = 8'b11000000;
    mem_c[1974] = 8'b11111111;
    mem_c[1975] = 8'b11111111;
    mem_c[1976] = 8'b11111111;
    mem_c[1977] = 8'b11111111;
    mem_c[1978] = 8'b11111111;
    mem_c[1979] = 8'b01111111;
    mem_c[1980] = 8'b00000000;
    mem_c[1981] = 8'b00000000;
    mem_c[1982] = 8'b00000000;
    mem_c[1983] = 8'b00000000;
    mem_c[1984] = 8'b00000000;
    mem_c[1985] = 8'b00000000;
    mem_c[1986] = 8'b00000000;
    mem_c[1987] = 8'b00000000;
    mem_c[1988] = 8'b00000000;
    mem_c[1989] = 8'b11000000;
    mem_c[1990] = 8'b11111111;
    mem_c[1991] = 8'b11111111;
    mem_c[1992] = 8'b11111111;
    mem_c[1993] = 8'b11111111;
    mem_c[1994] = 8'b11111111;
    mem_c[1995] = 8'b01111111;
    mem_c[1996] = 8'b00000000;
    mem_c[1997] = 8'b00000000;
    mem_c[1998] = 8'b00000000;
    mem_c[1999] = 8'b00000000;
    mem_c[2000] = 8'b00000000;
    mem_c[2001] = 8'b00000000;
    mem_c[2002] = 8'b00000000;
    mem_c[2003] = 8'b00000000;
    mem_c[2004] = 8'b00000000;
    mem_c[2005] = 8'b11000000;
    mem_c[2006] = 8'b11111111;
    mem_c[2007] = 8'b11111111;
    mem_c[2008] = 8'b11111111;
    mem_c[2009] = 8'b11111111;
    mem_c[2010] = 8'b11111111;
    mem_c[2011] = 8'b01111111;
    mem_c[2012] = 8'b00000000;
    mem_c[2013] = 8'b00000000;
    mem_c[2014] = 8'b00000000;
    mem_c[2015] = 8'b00000000;
    mem_c[2016] = 8'b00000000;
    mem_c[2017] = 8'b00000000;
    mem_c[2018] = 8'b00000000;
    mem_c[2019] = 8'b00000000;
    mem_c[2020] = 8'b00000000;
    mem_c[2021] = 8'b11000000;
    mem_c[2022] = 8'b11111111;
    mem_c[2023] = 8'b11111111;
    mem_c[2024] = 8'b11111111;
    mem_c[2025] = 8'b11111111;
    mem_c[2026] = 8'b11111111;
    mem_c[2027] = 8'b01111111;
    mem_c[2028] = 8'b00000000;
    mem_c[2029] = 8'b00000000;
    mem_c[2030] = 8'b00000000;
    mem_c[2031] = 8'b00000000;
    mem_c[2032] = 8'b00000000;
    mem_c[2033] = 8'b00000000;
    mem_c[2034] = 8'b00000000;
    mem_c[2035] = 8'b00000000;
    mem_c[2036] = 8'b00000000;
    mem_c[2037] = 8'b11111000;
    mem_c[2038] = 8'b11111111;
    mem_c[2039] = 8'b11111111;
    mem_c[2040] = 8'b11111111;
    mem_c[2041] = 8'b11111111;
    mem_c[2042] = 8'b11111111;
    mem_c[2043] = 8'b11111111;
    mem_c[2044] = 8'b00000011;
    mem_c[2045] = 8'b00000000;
    mem_c[2046] = 8'b00000000;
    mem_c[2047] = 8'b00000000;
end





  wire [10:0] addr = {y[6:0], x[6:3]};
  assign pixel = {mem_a[addr][x&7], mem_b[addr][x&7], mem_c[addr][x&7]};

endmodule
